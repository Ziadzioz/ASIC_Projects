module DLY1X1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX40M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX32M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX40M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX12M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module TIEHIM (
	Y, 
	VDD, 
	VSS);
   output Y;
   inout VDD;
   inout VSS;
endmodule

module TIELOM (
	Y, 
	VDD, 
	VSS);
   output Y;
   inout VDD;
   inout VSS;
endmodule

module BUFX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX5M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AO2B2X4M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AO2B2X2M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX2M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module NOR4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND4BX1M (
	Y, 
	D, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NAND3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI211X2M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFSQX2M (
	SN, 
	SI, 
	SE, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SN;
   input SI;
   input SE;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module MX2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AO2B2X1M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AND3X1M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKXOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI21BX1M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module XNOR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX1M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NOR4BX1M (
	Y, 
	D, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module CLKNAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MXI2X1M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module ADDHX1M (
	S, 
	CO, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module TLATNCAX12M (
	ECK, 
	E, 
	CK, 
	VDD, 
	VSS);
   output ECK;
   input E;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFQX2M (
	SI, 
	SE, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SEDFFX2M (
	SI, 
	SE, 
	QN, 
	Q, 
	E, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   output QN;
   output Q;
   input E;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module AO22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI31X1M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI32X1M (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI221XLM (
	Y, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI32X1M (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI31X2M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI21BX2M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OA21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1X1M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module NOR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AO21XLM (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX1M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OAI2B2X1M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module XNOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR3X1M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND4BBX1M (
	Y, 
	D, 
	C, 
	BN, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input BN;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AOI31X1M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX4M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB2X1M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module NOR3BX2M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module XOR3XLM (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND4X2M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI211X2M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module MX4X1M (
	Y, 
	S1, 
	S0, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S1;
   input S0;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI21BX1M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2B1X1M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND3BX2M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NAND3BX4M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module SDFFRX1M (
	SI, 
	SE, 
	RN, 
	QN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output QN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module OAI22X2M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI221X1M (
	Y, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1X2M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND4X2M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI222X1M (
	Y, 
	C1, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C1;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI222X1M (
	Y, 
	C1, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C1;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB2XLM (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module AOI21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI211X1M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI211X1M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OA21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2B11X1M (
	Y, 
	C0, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module ADDFX2M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKMX2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB1X1M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : K-2015.06
// Date      : Sat Aug 17 18:02:08 2024
/////////////////////////////////////////////////////////////
module DFT_MUX_0 (
	in_0, 
	in_1, 
	sel, 
	out, 
	VDD, 
	VSS);
   input in_0;
   input in_1;
   input sel;
   output out;
   inout VDD;
   inout VSS;

   // Module instantiations
   AO2B2X4M U1 (
	.Y(out),
	.B1(in_1),
	.B0(sel),
	.A1N(sel),
	.A0(in_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DFT_MUX_6 (
	in_0, 
	in_1, 
	sel, 
	out, 
	VDD, 
	VSS);
   input in_0;
   input in_1;
   input sel;
   output out;
   inout VDD;
   inout VSS;

   // Module instantiations
   AO2B2X4M U1 (
	.Y(out),
	.B1(in_1),
	.B0(sel),
	.A1N(sel),
	.A0(in_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DFT_MUX_5 (
	in_0, 
	in_1, 
	sel, 
	out, 
	VDD, 
	VSS);
   input in_0;
   input in_1;
   input sel;
   output out;
   inout VDD;
   inout VSS;

   // Module instantiations
   AO2B2X4M U1 (
	.Y(out),
	.B1(in_1),
	.B0(sel),
	.A1N(sel),
	.A0(in_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DFT_MUX_4 (
	in_0, 
	in_1, 
	sel, 
	out, 
	VDD, 
	VSS);
   input in_0;
   input in_1;
   input sel;
   output out;
   inout VDD;
   inout VSS;

   // Module instantiations
   AO2B2X4M U1 (
	.Y(out),
	.B1(in_1),
	.B0(sel),
	.A1N(sel),
	.A0(in_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DFT_MUX_3 (
	in_0, 
	in_1, 
	sel, 
	out, 
	VDD, 
	VSS);
   input in_0;
   input in_1;
   input sel;
   output out;
   inout VDD;
   inout VSS;

   // Module instantiations
   AO2B2X2M U1 (
	.Y(out),
	.B1(in_1),
	.B0(sel),
	.A1N(sel),
	.A0(in_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DFT_MUX_2 (
	in_0, 
	in_1, 
	sel, 
	out, 
	VDD, 
	VSS);
   input in_0;
   input in_1;
   input sel;
   output out;
   inout VDD;
   inout VSS;

   // Module instantiations
   AO2B2X4M U1 (
	.Y(out),
	.B1(in_1),
	.B0(sel),
	.A1N(sel),
	.A0(in_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DFT_MUX_1 (
	in_0, 
	in_1, 
	sel, 
	out, 
	VDD, 
	VSS);
   input in_0;
   input in_1;
   input sel;
   output out;
   inout VDD;
   inout VSS;

   // Module instantiations
   AO2B2X2M U1 (
	.Y(out),
	.B1(in_1),
	.B0(sel),
	.A1N(sel),
	.A0(in_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RESET_SYNC_NUM_STAGES2_test_0 (
	CLK, 
	RST, 
	RST_SYNC, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   output RST_SYNC;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire [1:0] SYNC_BUS;

   assign test_so = SYNC_BUS[1] ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M RST_SYNC_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(RST_SYNC),
	.D(SYNC_BUS[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[0]  (
	.SI(RST_SYNC),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_BUS[0]),
	.D(HTIE_LTIEHI_NET),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[1]  (
	.SI(SYNC_BUS[0]),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_BUS[1]),
	.D(SYNC_BUS[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RESET_SYNC_NUM_STAGES2_test_1 (
	CLK, 
	RST, 
	RST_SYNC, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   output RST_SYNC;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire [1:0] SYNC_BUS;

   assign test_so = SYNC_BUS[1] ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M RST_SYNC_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(RST_SYNC),
	.D(SYNC_BUS[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[0]  (
	.SI(RST_SYNC),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_BUS[0]),
	.D(HTIE_LTIEHI_NET),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[1]  (
	.SI(SYNC_BUS[0]),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_BUS[1]),
	.D(SYNC_BUS[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module PRESCALE_BLOCK (
	PRESCALE, 
	DIV_RATIO, 
	VDD, 
	VSS);
   input [5:0] PRESCALE;
   output [7:0] DIV_RATIO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n1;
   wire n2;
   wire n3;
   wire n4;

   assign DIV_RATIO[4] = 1'b0 ;
   assign DIV_RATIO[5] = 1'b0 ;
   assign DIV_RATIO[6] = 1'b0 ;
   assign DIV_RATIO[7] = 1'b0 ;

   // Module instantiations
   NOR4X1M U3 (
	.Y(DIV_RATIO[3]),
	.D(PRESCALE[4]),
	.C(PRESCALE[5]),
	.B(PRESCALE[3]),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U4 (
	.Y(DIV_RATIO[2]),
	.C(PRESCALE[0]),
	.B(PRESCALE[1]),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U5 (
	.Y(n6),
	.D(n1),
	.C(n2),
	.B(PRESCALE[3]),
	.AN(PRESCALE[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U6 (
	.Y(n7),
	.D(n1),
	.C(n2),
	.B(PRESCALE[4]),
	.AN(PRESCALE[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U7 (
	.Y(DIV_RATIO[1]),
	.C(PRESCALE[0]),
	.B(PRESCALE[1]),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U8 (
	.Y(n5),
	.C(PRESCALE[2]),
	.B(n3),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U9 (
	.Y(DIV_RATIO[0]),
	.C0(n3),
	.B0(n4),
	.A1(n9),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U10 (
	.Y(n9),
	.B(n6),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U11 (
	.Y(n8),
	.D(n2),
	.C(PRESCALE[3]),
	.B(PRESCALE[4]),
	.A(PRESCALE[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(n3),
	.A(PRESCALE[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U13 (
	.Y(n2),
	.A(PRESCALE[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U14 (
	.Y(n4),
	.A(PRESCALE[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U15 (
	.Y(n1),
	.A(PRESCALE[5]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module CLK_DIV_test_1 (
	RST_EN, 
	I_REF_CLK, 
	CLK_EN, 
	DIV_RATIO, 
	O_DIV_CLK, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN0_scanrst1, 
	n12__Exclude_0_NET, 
	scanclkuart__L4_N0, 
	scanclkuart__L6_N0, 
	VDD, 
	VSS);
   input RST_EN;
   input I_REF_CLK;
   input CLK_EN;
   input [7:0] DIV_RATIO;
   output O_DIV_CLK;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN0_scanrst1;
   input n12__Exclude_0_NET;
   input scanclkuart__L4_N0;
   input scanclkuart__L6_N0;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire out_clk;
   wire flag;
   wire N13;
   wire N14;
   wire N15;
   wire N16;
   wire N17;
   wire N18;
   wire N19;
   wire N20;
   wire N25;
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire N32;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire [7:0] counter;

//   assign test_so = out_clk ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M flag_reg (
	.SN(RST_EN),
	.SI(counter[7]),
	.SE(test_se),
	.Q(flag),
	.D(n29),
	.CK(scanclkuart__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M out_clk_reg (
	.SI(flag),
	.SE(test_se),
	.RN(RST_EN),
	.Q(test_so),
	.D(n30),
	.CK(I_REF_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[7]  (
	.SI(counter[6]),
	.SE(test_se),
	.RN(FE_OFN0_scanrst1),
	.Q(counter[7]),
	.D(n31),
	.CK(scanclkuart__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(FE_OFN0_scanrst1),
	.Q(counter[0]),
	.D(n38),
	.CK(scanclkuart__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[6]  (
	.SI(counter[5]),
	.SE(test_se),
	.RN(FE_OFN0_scanrst1),
	.Q(counter[6]),
	.D(n32),
	.CK(scanclkuart__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[5]  (
	.SI(counter[4]),
	.SE(test_se),
	.RN(FE_OFN0_scanrst1),
	.Q(counter[5]),
	.D(n33),
	.CK(scanclkuart__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[4]  (
	.SI(counter[3]),
	.SE(test_se),
	.RN(FE_OFN0_scanrst1),
	.Q(counter[4]),
	.D(n34),
	.CK(scanclkuart__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[3]  (
	.SI(counter[2]),
	.SE(test_se),
	.RN(FE_OFN0_scanrst1),
	.Q(counter[3]),
	.D(n35),
	.CK(scanclkuart__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[2]  (
	.SI(counter[1]),
	.SE(test_se),
	.RN(RST_EN),
	.Q(counter[2]),
	.D(n36),
	.CK(scanclkuart__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[1]  (
	.SI(counter[0]),
	.SE(test_se),
	.RN(RST_EN),
	.Q(counter[1]),
	.D(n37),
	.CK(scanclkuart__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U5 (
	.Y(n51),
	.B(n18),
	.AN(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U7 (
	.Y(O_DIV_CLK),
	.S0(n51),
	.B(test_so),
	.A(scanclkuart__L4_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X1M U12 (
	.Y(n38),
	.B1(n1),
	.B0(N25),
	.A1N(n51),
	.A0(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X1M U17 (
	.Y(n37),
	.B1(n1),
	.B0(N26),
	.A1N(n51),
	.A0(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X1M U18 (
	.Y(n36),
	.B1(n1),
	.B0(N27),
	.A1N(n51),
	.A0(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X1M U19 (
	.Y(n35),
	.B1(n1),
	.B0(N28),
	.A1N(n51),
	.A0(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X1M U20 (
	.Y(n34),
	.B1(n1),
	.B0(N29),
	.A1N(n51),
	.A0(counter[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X1M U21 (
	.Y(n33),
	.B1(n1),
	.B0(N30),
	.A1N(n51),
	.A0(counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X1M U22 (
	.Y(n32),
	.B1(n1),
	.B0(N31),
	.A1N(n51),
	.A0(counter[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X1M U23 (
	.Y(n31),
	.B1(n1),
	.B0(N32),
	.A1N(n51),
	.A0(counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X1M U24 (
	.Y(n1),
	.C(n51),
	.B(n4),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U25 (
	.Y(n30),
	.B(n5),
	.A(n12__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21BX1M U26 (
	.Y(n5),
	.B0N(n51),
	.A1(n3),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U27 (
	.Y(n3),
	.B(DIV_RATIO[0]),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U28 (
	.Y(n29),
	.B(n7),
	.A(flag), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U29 (
	.Y(n7),
	.B(n51),
	.AN(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4BX1M U30 (
	.Y(n18),
	.D(DIV_RATIO[1]),
	.C(DIV_RATIO[3]),
	.B(DIV_RATIO[2]),
	.AN(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U31 (
	.Y(n19),
	.D(DIV_RATIO[4]),
	.C(DIV_RATIO[5]),
	.B(DIV_RATIO[6]),
	.A(DIV_RATIO[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U32 (
	.Y(n4),
	.B(DIV_RATIO[0]),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U33 (
	.Y(n20),
	.S0(flag),
	.B(n6),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U34 (
	.Y(n6),
	.B(n23),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U35 (
	.Y(n23),
	.D(n26),
	.C(n25),
	.B(n24),
	.A(counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U36 (
	.Y(n26),
	.B(DIV_RATIO[3]),
	.A(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U37 (
	.Y(n25),
	.B(DIV_RATIO[2]),
	.A(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U38 (
	.Y(n24),
	.B(DIV_RATIO[1]),
	.A(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U39 (
	.Y(n22),
	.D(n40),
	.C(n39),
	.B(n28),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U40 (
	.Y(n40),
	.B(DIV_RATIO[7]),
	.A(counter[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U41 (
	.Y(n39),
	.B(DIV_RATIO[6]),
	.A(counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U42 (
	.Y(n28),
	.B(DIV_RATIO[5]),
	.A(counter[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U43 (
	.Y(n27),
	.B(DIV_RATIO[4]),
	.A(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U44 (
	.Y(n21),
	.B(n42),
	.A(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U45 (
	.Y(n42),
	.D(n46),
	.C(n45),
	.B(n44),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U46 (
	.Y(n46),
	.B(N16),
	.A(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U47 (
	.Y(n45),
	.B(N15),
	.A(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U48 (
	.Y(n44),
	.B(N14),
	.A(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U49 (
	.Y(n43),
	.B(N13),
	.A(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U50 (
	.Y(n41),
	.D(n50),
	.C(n49),
	.B(n48),
	.A(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U51 (
	.Y(n50),
	.B(N20),
	.A(counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U52 (
	.Y(n49),
	.B(N19),
	.A(counter[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U53 (
	.Y(n48),
	.B(N18),
	.A(counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U54 (
	.Y(n47),
	.B(N17),
	.A(counter[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLK_DIV_0_DW01_inc_0 add_43 (
	.A({ counter[7],
		counter[6],
		counter[5],
		counter[4],
		counter[3],
		counter[2],
		counter[1],
		counter[0] }),
	.SUM({ N32,
		N31,
		N30,
		N29,
		N28,
		N27,
		N26,
		N25 }), 
	.VDD(VDD), 
	.VSS(VSS));
   CLK_DIV_0_DW01_inc_1 add_36 (
	.A({ 1'b0,
		DIV_RATIO[7],
		DIV_RATIO[6],
		DIV_RATIO[5],
		DIV_RATIO[4],
		DIV_RATIO[3],
		DIV_RATIO[2],
		DIV_RATIO[1] }),
	.SUM({ N20,
		N19,
		N18,
		N17,
		N16,
		N15,
		N14,
		N13 }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module CLK_DIV_0_DW01_inc_0 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [7:0] A;
   output [7:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [7:2] carry;

   // Module instantiations
   ADDHX1M U1_1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.B(carry[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U1 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U2 (
	.Y(SUM[7]),
	.B(A[7]),
	.A(carry[7]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module CLK_DIV_0_DW01_inc_1 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [7:0] A;
   output [7:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [7:2] carry;

   // Module instantiations
   ADDHX1M U1_1_6 (
	.S(SUM[6]),
	.CO(SUM[7]),
	.B(carry[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U1 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module CLK_DIV_test_0 (
	RST_EN, 
	I_REF_CLK, 
	CLK_EN, 
	DIV_RATIO, 
	O_DIV_CLK, 
	test_si, 
	test_so, 
	test_se, 
	n13__Exclude_0_NET, 
	scanclkuart__L4_N0, 
	scanclkuart__L6_N0, 
	VDD, 
	VSS);
   input RST_EN;
   input I_REF_CLK;
   input CLK_EN;
   input [7:0] DIV_RATIO;
   output O_DIV_CLK;
   input test_si;
   output test_so;
   input test_se;
   input n13__Exclude_0_NET;
   input scanclkuart__L4_N0;
   input scanclkuart__L6_N0;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire LTIE_LTIELO_NET;
   wire out_clk;
   wire flag;
   wire N13;
   wire N14;
   wire N15;
   wire N16;
   wire N17;
   wire N18;
   wire N19;
   wire N20;
   wire N25;
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire N32;
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire [7:0] counter;

//   assign test_so = out_clk ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M flag_reg (
	.SN(RST_EN),
	.SI(counter[7]),
	.SE(test_se),
	.Q(flag),
	.D(n61),
	.CK(scanclkuart__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M out_clk_reg (
	.SI(flag),
	.SE(test_se),
	.RN(RST_EN),
	.Q(test_so),
	.D(n60),
	.CK(I_REF_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[7]  (
	.SI(counter[6]),
	.SE(test_se),
	.RN(RST_EN),
	.Q(counter[7]),
	.D(n59),
	.CK(scanclkuart__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST_EN),
	.Q(counter[0]),
	.D(n52),
	.CK(scanclkuart__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[6]  (
	.SI(counter[5]),
	.SE(test_se),
	.RN(RST_EN),
	.Q(counter[6]),
	.D(n58),
	.CK(scanclkuart__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[5]  (
	.SI(counter[4]),
	.SE(test_se),
	.RN(RST_EN),
	.Q(counter[5]),
	.D(n57),
	.CK(scanclkuart__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[4]  (
	.SI(counter[3]),
	.SE(test_se),
	.RN(RST_EN),
	.Q(counter[4]),
	.D(n56),
	.CK(scanclkuart__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[3]  (
	.SI(counter[2]),
	.SE(test_se),
	.RN(RST_EN),
	.Q(counter[3]),
	.D(n55),
	.CK(scanclkuart__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[2]  (
	.SI(counter[1]),
	.SE(test_se),
	.RN(RST_EN),
	.Q(counter[2]),
	.D(n54),
	.CK(scanclkuart__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[1]  (
	.SI(counter[0]),
	.SE(test_se),
	.RN(RST_EN),
	.Q(counter[1]),
	.D(n53),
	.CK(scanclkuart__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U5 (
	.Y(n51),
	.B(n18),
	.AN(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U7 (
	.Y(O_DIV_CLK),
	.S0(n51),
	.B(test_so),
	.A(scanclkuart__L4_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X1M U12 (
	.Y(n52),
	.B1(n1),
	.B0(N25),
	.A1N(n51),
	.A0(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X1M U17 (
	.Y(n53),
	.B1(n1),
	.B0(N26),
	.A1N(n51),
	.A0(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X1M U18 (
	.Y(n54),
	.B1(n1),
	.B0(N27),
	.A1N(n51),
	.A0(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X1M U19 (
	.Y(n55),
	.B1(n1),
	.B0(N28),
	.A1N(n51),
	.A0(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X1M U20 (
	.Y(n56),
	.B1(n1),
	.B0(N29),
	.A1N(n51),
	.A0(counter[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X1M U21 (
	.Y(n57),
	.B1(n1),
	.B0(N30),
	.A1N(n51),
	.A0(counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X1M U22 (
	.Y(n58),
	.B1(n1),
	.B0(N31),
	.A1N(n51),
	.A0(counter[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X1M U23 (
	.Y(n59),
	.B1(n1),
	.B0(N32),
	.A1N(n51),
	.A0(counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X1M U24 (
	.Y(n1),
	.C(n51),
	.B(n4),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U25 (
	.Y(n60),
	.B(n5),
	.A(n13__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21BX1M U26 (
	.Y(n5),
	.B0N(n51),
	.A1(n3),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U27 (
	.Y(n3),
	.B(DIV_RATIO[0]),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U28 (
	.Y(n61),
	.B(n7),
	.A(flag), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U29 (
	.Y(n7),
	.B(n51),
	.AN(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4BX1M U30 (
	.Y(n18),
	.D(DIV_RATIO[1]),
	.C(DIV_RATIO[3]),
	.B(DIV_RATIO[2]),
	.AN(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U31 (
	.Y(n19),
	.D(LTIE_LTIELO_NET),
	.C(LTIE_LTIELO_NET),
	.B(LTIE_LTIELO_NET),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U32 (
	.Y(n4),
	.B(DIV_RATIO[0]),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U33 (
	.Y(n20),
	.S0(flag),
	.B(n6),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U34 (
	.Y(n6),
	.B(n23),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U35 (
	.Y(n23),
	.D(n26),
	.C(n25),
	.B(n24),
	.A(counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U36 (
	.Y(n26),
	.B(DIV_RATIO[3]),
	.A(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U37 (
	.Y(n25),
	.B(DIV_RATIO[2]),
	.A(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U38 (
	.Y(n24),
	.B(DIV_RATIO[1]),
	.A(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U39 (
	.Y(n22),
	.D(n40),
	.C(n39),
	.B(n28),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U40 (
	.Y(n40),
	.B(LTIE_LTIELO_NET),
	.A(counter[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U41 (
	.Y(n39),
	.B(LTIE_LTIELO_NET),
	.A(counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U42 (
	.Y(n28),
	.B(LTIE_LTIELO_NET),
	.A(counter[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U43 (
	.Y(n27),
	.B(LTIE_LTIELO_NET),
	.A(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U44 (
	.Y(n21),
	.B(n42),
	.A(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U45 (
	.Y(n42),
	.D(n46),
	.C(n45),
	.B(n44),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U46 (
	.Y(n46),
	.B(N16),
	.A(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U47 (
	.Y(n45),
	.B(N15),
	.A(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U48 (
	.Y(n44),
	.B(N14),
	.A(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U49 (
	.Y(n43),
	.B(N13),
	.A(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U50 (
	.Y(n41),
	.D(n50),
	.C(n49),
	.B(n48),
	.A(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U51 (
	.Y(n50),
	.B(N20),
	.A(counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U52 (
	.Y(n49),
	.B(N19),
	.A(counter[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U53 (
	.Y(n48),
	.B(N18),
	.A(counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U54 (
	.Y(n47),
	.B(N17),
	.A(counter[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLK_DIV_1_DW01_inc_0 add_43 (
	.A({ counter[7],
		counter[6],
		counter[5],
		counter[4],
		counter[3],
		counter[2],
		counter[1],
		counter[0] }),
	.SUM({ N32,
		N31,
		N30,
		N29,
		N28,
		N27,
		N26,
		N25 }), 
	.VDD(VDD), 
	.VSS(VSS));
   CLK_DIV_1_DW01_inc_1 add_36 (
	.A({ 1'b0,
		DIV_RATIO[7],
		DIV_RATIO[6],
		DIV_RATIO[5],
		DIV_RATIO[4],
		DIV_RATIO[3],
		DIV_RATIO[2],
		DIV_RATIO[1] }),
	.SUM({ N20,
		N19,
		N18,
		N17,
		N16,
		N15,
		N14,
		N13 }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module CLK_DIV_1_DW01_inc_0 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [7:0] A;
   output [7:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [7:2] carry;

   // Module instantiations
   ADDHX1M U1_1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.B(carry[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U1 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U2 (
	.Y(SUM[7]),
	.B(A[7]),
	.A(carry[7]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module CLK_DIV_1_DW01_inc_1 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [7:0] A;
   output [7:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire LTIE_LTIELO_NET;
   wire [7:2] carry;

   // Module instantiations
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_6 (
	.S(SUM[6]),
	.CO(SUM[7]),
	.B(carry[6]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U1 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module CLOCK_GATING (
	REF_CLK, 
	CLK_GATE_EN, 
	ALU_CLK, 
	VDD, 
	VSS);
   input REF_CLK;
   input CLK_GATE_EN;
   output ALU_CLK;
   inout VDD;
   inout VSS;

   // Module instantiations
   TLATNCAX12M U0_TLATNCAX12M (
	.ECK(ALU_CLK),
	.E(CLK_GATE_EN),
	.CK(REF_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module PULSE_GENRATOR_BLOCK_test_1 (
	TX_CLK, 
	PULSE_GEN, 
	RINC, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input TX_CLK;
   input PULSE_GEN;
   output RINC;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire BEFORE_INV;
   wire AFTER_INV;

   // Module instantiations
   SDFFQX2M BEFORE_INV_reg (
	.SI(test_si),
	.SE(test_se),
	.Q(BEFORE_INV),
	.D(PULSE_GEN),
	.CK(TX_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M RINC_reg (
	.SI(BEFORE_INV),
	.SE(test_se),
	.Q(RINC),
	.D(AFTER_INV),
	.CK(TX_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U5 (
	.Y(AFTER_INV),
	.B(BEFORE_INV),
	.AN(PULSE_GEN), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DATA_SYNC_NUM_STAGES2_BUS_WIDTH8_test_1 (
	CLK, 
	RST, 
	EN, 
	UNSYNC_BUS, 
	enable_pulse, 
	SYNC_BUS, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN1_scanrst2, 
	FE_OFN3_scanclkref, 
	FE_OFN11_SE, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input EN;
   input [7:0] UNSYNC_BUS;
   output enable_pulse;
   output [7:0] SYNC_BUS;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN1_scanrst2;
   input FE_OFN3_scanclkref;
   input FE_OFN11_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n2;
   wire n4;
   wire n6;
   wire n8;
   wire n10;
   wire n12;
   wire n14;
   wire n16;
   wire n18;
   wire n23;
   wire [1:0] bus_en_sync;

   // Module instantiations
   SEDFFX2M pulse_reg (
	.SI(enable_pulse),
	.SE(FE_OFN11_SE),
	.QN(n2),
	.Q(test_so),
	.E(RST),
	.D(bus_en_sync[1]),
	.CK(FE_OFN3_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SEDFFX2M \bus_en_sync_reg[1]  (
	.SI(bus_en_sync[0]),
	.SE(FE_OFN11_SE),
	.Q(bus_en_sync[1]),
	.E(RST),
	.D(bus_en_sync[0]),
	.CK(FE_OFN3_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[7]  (
	.SI(SYNC_BUS[6]),
	.SE(test_se),
	.RN(FE_OFN1_scanrst2),
	.Q(SYNC_BUS[7]),
	.D(n18),
	.CK(FE_OFN3_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[4]  (
	.SI(SYNC_BUS[3]),
	.SE(test_se),
	.RN(FE_OFN1_scanrst2),
	.Q(SYNC_BUS[4]),
	.D(n12),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[3]  (
	.SI(SYNC_BUS[2]),
	.SE(test_se),
	.RN(FE_OFN1_scanrst2),
	.Q(SYNC_BUS[3]),
	.D(n10),
	.CK(FE_OFN3_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[1]  (
	.SI(SYNC_BUS[0]),
	.SE(test_se),
	.RN(FE_OFN1_scanrst2),
	.Q(SYNC_BUS[1]),
	.D(n6),
	.CK(FE_OFN3_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[5]  (
	.SI(SYNC_BUS[4]),
	.SE(test_se),
	.RN(FE_OFN1_scanrst2),
	.Q(SYNC_BUS[5]),
	.D(n14),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[0]  (
	.SI(test_si),
	.SE(FE_OFN11_SE),
	.RN(RST),
	.Q(SYNC_BUS[0]),
	.D(n4),
	.CK(FE_OFN3_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[2]  (
	.SI(SYNC_BUS[1]),
	.SE(test_se),
	.RN(FE_OFN1_scanrst2),
	.Q(SYNC_BUS[2]),
	.D(n8),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[6]  (
	.SI(SYNC_BUS[5]),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_BUS[6]),
	.D(n16),
	.CK(FE_OFN3_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M enable_pulse_reg (
	.SI(bus_en_sync[1]),
	.SE(FE_OFN11_SE),
	.RN(RST),
	.Q(enable_pulse),
	.D(n23),
	.CK(FE_OFN3_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SEDFFX2M \bus_en_sync_reg[0]  (
	.SI(SYNC_BUS[7]),
	.SE(test_se),
	.Q(bus_en_sync[0]),
	.E(FE_OFN1_scanrst2),
	.D(EN),
	.CK(FE_OFN3_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(n23),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U4 (
	.Y(n1),
	.B(n2),
	.A(bus_en_sync[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U5 (
	.Y(n4),
	.B1(n1),
	.B0(SYNC_BUS[0]),
	.A1(n23),
	.A0(UNSYNC_BUS[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U6 (
	.Y(n6),
	.B1(n1),
	.B0(SYNC_BUS[1]),
	.A1(n23),
	.A0(UNSYNC_BUS[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U7 (
	.Y(n8),
	.B1(n1),
	.B0(SYNC_BUS[2]),
	.A1(n23),
	.A0(UNSYNC_BUS[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U8 (
	.Y(n10),
	.B1(n1),
	.B0(SYNC_BUS[3]),
	.A1(n23),
	.A0(UNSYNC_BUS[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U9 (
	.Y(n12),
	.B1(n1),
	.B0(SYNC_BUS[4]),
	.A1(n23),
	.A0(UNSYNC_BUS[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U10 (
	.Y(n14),
	.B1(n1),
	.B0(SYNC_BUS[5]),
	.A1(n23),
	.A0(UNSYNC_BUS[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U11 (
	.Y(n16),
	.B1(n1),
	.B0(SYNC_BUS[6]),
	.A1(n23),
	.A0(UNSYNC_BUS[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U12 (
	.Y(n18),
	.B1(n1),
	.B0(SYNC_BUS[7]),
	.A1(n23),
	.A0(UNSYNC_BUS[7]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SYS_UART_TOP_DATA_WIDTH8_test_1 (
	TX_CLK, 
	RX_CLK, 
	RST_SYNC_1, 
	RX_IN, 
	R_EMPTY, 
	UART_CONFIG, 
	R_DATA, 
	Tx_OUT, 
	DATA_VALID, 
	Stop_error, 
	Parity_error, 
	PULSE_GEN, 
	P_DATA, 
	test_si, 
	test_se, 
	FE_OFN0_scanrst1, 
	FE_OFN11_SE, 
	FE_OFN12_SE, 
	FE_OFN13_SE, 
	FE_OFN14_SE, 
	VDD, 
	VSS);
   input TX_CLK;
   input RX_CLK;
   input RST_SYNC_1;
   input RX_IN;
   input R_EMPTY;
   input [7:0] UART_CONFIG;
   input [7:0] R_DATA;
   output Tx_OUT;
   output DATA_VALID;
   output Stop_error;
   output Parity_error;
   output PULSE_GEN;
   output [7:0] P_DATA;
   input test_si;
   input test_se;
   input FE_OFN0_scanrst1;
   input FE_OFN11_SE;
   input FE_OFN12_SE;
   input FE_OFN13_SE;
   input FE_OFN14_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n2;
   wire n3;

   // Module instantiations
   UART_RX_TOP_test_1 UART_RX_TOP (
	.CLK(RX_CLK),
	.RST(RST_SYNC_1),
	.RX_IN(RX_IN),
	.Parity_en(UART_CONFIG[0]),
	.Parity_type(UART_CONFIG[1]),
	.Prescale({ UART_CONFIG[7],
		UART_CONFIG[6],
		UART_CONFIG[5],
		UART_CONFIG[4],
		UART_CONFIG[3],
		UART_CONFIG[2] }),
	.DATA_VALID(DATA_VALID),
	.Stop_error(Stop_error),
	.Parity_error(Parity_error),
	.P_DATA({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }),
	.test_si2(n2),
	.test_si1(test_si),
	.test_so1(n3),
	.test_se(test_se),
	.FE_OFN0_scanrst1(FE_OFN0_scanrst1),
	.FE_OFN11_SE(FE_OFN11_SE),
	.FE_OFN14_SE(FE_OFN14_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   UART_TX_TOP_DATA_WIDTH8_test_1 UART_TX_TOP (
	.CLK(TX_CLK),
	.RST(FE_OFN0_scanrst1),
	.party_en(UART_CONFIG[0]),
	.data_valid(R_EMPTY),
	.party_typ(UART_CONFIG[1]),
	.P_DATA({ R_DATA[7],
		R_DATA[6],
		R_DATA[5],
		R_DATA[4],
		R_DATA[3],
		R_DATA[2],
		R_DATA[1],
		R_DATA[0] }),
	.busy(PULSE_GEN),
	.Tx_OUT(Tx_OUT),
	.test_si(n3),
	.test_so(n2),
	.test_se(FE_OFN12_SE),
	.FE_OFN13_SE(FE_OFN13_SE), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_RX_TOP_test_1 (
	CLK, 
	RST, 
	RX_IN, 
	Parity_en, 
	Parity_type, 
	Prescale, 
	DATA_VALID, 
	Stop_error, 
	Parity_error, 
	P_DATA, 
	test_si2, 
	test_si1, 
	test_so1, 
	test_se, 
	FE_OFN0_scanrst1, 
	FE_OFN11_SE, 
	FE_OFN14_SE, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input RX_IN;
   input Parity_en;
   input Parity_type;
   input [5:0] Prescale;
   output DATA_VALID;
   output Stop_error;
   output Parity_error;
   output [7:0] P_DATA;
   input test_si2;
   input test_si1;
   output test_so1;
   input test_se;
   input FE_OFN0_scanrst1;
   input FE_OFN11_SE;
   input FE_OFN14_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire Start_glitch;
   wire Data_samp_en;
   wire edge_count_en;
   wire desrializer_en;
   wire stop_en;
   wire start_en;
   wire parity_check_en;
   wire Sampled_Bit;
   wire parity_flag;
   wire n3;
   wire n4;
   wire [3:0] bit_count;
   wire [5:0] edge_count;

   assign test_so1 = Start_glitch ;

   // Module instantiations
   FSM_test_1 FSM (
	.CLK(CLK),
	.RST(RST),
	.RX_IN(RX_IN),
	.Parity_error(Parity_error),
	.Stop_error(Stop_error),
	.Start_glitch(Start_glitch),
	.Parity_en(Parity_en),
	.bit_count({ bit_count[3],
		bit_count[2],
		bit_count[1],
		bit_count[0] }),
	.edge_count({ edge_count[5],
		edge_count[4],
		edge_count[3],
		edge_count[2],
		edge_count[1],
		edge_count[0] }),
	.Data_samp_en(Data_samp_en),
	.edge_count_en(edge_count_en),
	.desrializer_en(desrializer_en),
	.stop_en(stop_en),
	.start_en(start_en),
	.parity_check_en(parity_check_en),
	.DATA_VALID(DATA_VALID),
	.test_si(parity_flag),
	.test_so(n3),
	.test_se(FE_OFN14_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   Bit_counter_test_1 Bit_counter (
	.CLK(CLK),
	.RST(RST),
	.edge_count_en(edge_count_en),
	.Prescale({ Prescale[5],
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }),
	.bit_count({ bit_count[3],
		bit_count[2],
		bit_count[1],
		bit_count[0] }),
	.edge_count({ edge_count[5],
		edge_count[4],
		edge_count[3],
		edge_count[2],
		edge_count[1],
		edge_count[0] }),
	.test_si(test_si1),
	.test_se(test_se),
	.FE_OFN14_SE(FE_OFN14_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   Data_Sampling_test_1 Data_Sampling (
	.CLK(CLK),
	.RST(RST),
	.Data_samp_en(Data_samp_en),
	.RX_IN(RX_IN),
	.Prescale({ Prescale[5],
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }),
	.edge_count({ edge_count[5],
		edge_count[4],
		edge_count[3],
		edge_count[2],
		edge_count[1],
		edge_count[0] }),
	.Sampled_Bit(Sampled_Bit),
	.test_so(n4),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   Start_Check_test_1 Start_Check (
	.CLK(CLK),
	.RST(FE_OFN0_scanrst1),
	.start_en(start_en),
	.Sampled_Bit(Sampled_Bit),
	.Start_glitch(Start_glitch),
	.test_si(Parity_error),
	.test_se(FE_OFN11_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   Stop_Check_test_1 Stop_Check (
	.CLK(CLK),
	.RST(FE_OFN0_scanrst1),
	.stop_en(stop_en),
	.Sampled_Bit(Sampled_Bit),
	.Stop_error(Stop_error),
	.test_si(test_si2),
	.test_se(FE_OFN14_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   Deserializer_test_1 Deserializer (
	.CLK(CLK),
	.RST(RST),
	.desrializer_en(desrializer_en),
	.Sampled_Bit(Sampled_Bit),
	.DATA_VALID(DATA_VALID),
	.bit_count({ bit_count[3],
		bit_count[2],
		bit_count[1],
		bit_count[0] }),
	.parity_flag(parity_flag),
	.P_DATA({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }),
	.test_si(n4),
	.test_se(test_se),
	.FE_OFN11_SE(FE_OFN11_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   Parity_Check_test_1 Parity_Check (
	.CLK(CLK),
	.RST(FE_OFN0_scanrst1),
	.Parity_type(Parity_type),
	.parity_check_en(parity_check_en),
	.Sampled_Bit(Sampled_Bit),
	.parity_flag(parity_flag),
	.Parity_error(Parity_error),
	.test_si(n3),
	.test_se(FE_OFN11_SE), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FSM_test_1 (
	CLK, 
	RST, 
	RX_IN, 
	Parity_error, 
	Stop_error, 
	Start_glitch, 
	Parity_en, 
	bit_count, 
	edge_count, 
	Data_samp_en, 
	edge_count_en, 
	desrializer_en, 
	stop_en, 
	start_en, 
	parity_check_en, 
	DATA_VALID, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input RX_IN;
   input Parity_error;
   input Stop_error;
   input Start_glitch;
   input Parity_en;
   input [3:0] bit_count;
   input [5:0] edge_count;
   output Data_samp_en;
   output edge_count_en;
   output desrializer_en;
   output stop_en;
   output start_en;
   output parity_check_en;
   output DATA_VALID;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n14;
   wire n15;
   wire n16;
   wire [2:0] current_state;
   wire [2:0] next_state;

   assign edge_count_en = Data_samp_en ;
   assign test_so = current_state[2] ;

   // Module instantiations
   SDFFRQX2M \current_state_reg[1]  (
	.SI(current_state[0]),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[1]),
	.D(next_state[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[0]),
	.D(next_state[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[2]  (
	.SI(current_state[1]),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[2]),
	.D(next_state[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U6 (
	.Y(n7),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U7 (
	.Y(DATA_VALID),
	.B(stop_en),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U8 (
	.Y(n22),
	.B(n8),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U9 (
	.Y(n26),
	.B(n22),
	.A(parity_check_en), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U10 (
	.Y(n14),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U11 (
	.Y(desrializer_en),
	.B0(n14),
	.A1(n37),
	.A0(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(n6),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U13 (
	.Y(Data_samp_en),
	.B0(stop_en),
	.A1(n38),
	.A0(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U14 (
	.Y(n40),
	.C(n11),
	.B(bit_count[2]),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U15 (
	.Y(parity_check_en),
	.C(n15),
	.B(current_state[2]),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U16 (
	.Y(n20),
	.C(n15),
	.B(current_state[2]),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U17 (
	.Y(n28),
	.C(n8),
	.B(bit_count[2]),
	.A(bit_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U18 (
	.Y(start_en),
	.C(n12),
	.B(current_state[2]),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U19 (
	.Y(next_state[2]),
	.B0(n19),
	.A2(n18),
	.A1(n4),
	.A0(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n4),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U21 (
	.Y(n19),
	.B1(parity_check_en),
	.B0(n21),
	.A2(n20),
	.A1(n16),
	.A0(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U22 (
	.Y(n18),
	.C0(n5),
	.B1(n16),
	.B0(n22),
	.A1(n23),
	.A0(Parity_en), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U23 (
	.Y(n24),
	.B(n5),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U24 (
	.Y(n33),
	.B1(n23),
	.B0(Parity_en),
	.A2(n10),
	.A1(n16),
	.A0(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U25 (
	.Y(n10),
	.A(bit_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U26 (
	.Y(n34),
	.C(bit_count[3]),
	.B(n9),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U27 (
	.Y(n38),
	.B(current_state[1]),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U28 (
	.Y(next_state[1]),
	.C0(n27),
	.B0(n26),
	.A1(n14),
	.A0(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U29 (
	.Y(n25),
	.B(n29),
	.A(Parity_en), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U30 (
	.Y(n27),
	.D(n28),
	.C(start_en),
	.B(n11),
	.AN(Start_glitch), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U31 (
	.Y(n8),
	.A(bit_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U32 (
	.Y(n23),
	.B(n40),
	.A(bit_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U33 (
	.Y(stop_en),
	.B(current_state[2]),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U34 (
	.Y(n29),
	.B(bit_count[3]),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U36 (
	.Y(n37),
	.B(n5),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U37 (
	.Y(n39),
	.B1(n23),
	.B0(n16),
	.A1(n22),
	.A0(Parity_en), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U38 (
	.Y(n9),
	.A(bit_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U39 (
	.Y(n5),
	.A(Stop_error), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U40 (
	.Y(n32),
	.B0(RX_IN),
	.A1(n24),
	.A0(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U41 (
	.Y(n17),
	.C(current_state[2]),
	.B(n15),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U42 (
	.Y(n15),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U43 (
	.Y(n12),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U44 (
	.Y(n21),
	.B(n22),
	.A(Parity_error), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U45 (
	.Y(n11),
	.A(bit_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U46 (
	.Y(next_state[0]),
	.B(n31),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U47 (
	.Y(n30),
	.B0(n35),
	.A2(Parity_en),
	.A1(n6),
	.A0(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U48 (
	.Y(n31),
	.B0(n7),
	.A2(n32),
	.A1(n15),
	.A0(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21BX2M U49 (
	.Y(n35),
	.B0N(start_en),
	.A1(n11),
	.A0(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U50 (
	.Y(n16),
	.A(Parity_en), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Bit_counter_test_1 (
	CLK, 
	RST, 
	edge_count_en, 
	Prescale, 
	bit_count, 
	edge_count, 
	test_si, 
	test_se, 
	FE_OFN14_SE, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input edge_count_en;
   input [5:0] Prescale;
   output [3:0] bit_count;
   output [5:0] edge_count;
   input test_si;
   input test_se;
   input FE_OFN14_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N7;
   wire N8;
   wire N9;
   wire N10;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire N20;
   wire N21;
   wire N22;
   wire N23;
   wire N24;
   wire N25;
   wire N36;
   wire N37;
   wire N38;
   wire N39;
   wire N40;
   wire N41;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire \add_27/carry[5] ;
   wire \add_27/carry[4] ;
   wire \add_27/carry[3] ;
   wire \add_27/carry[2] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;

   // Module instantiations
   SDFFRQX2M \edge_count_reg[5]  (
	.SI(edge_count[4]),
	.SE(test_se),
	.RN(RST),
	.Q(edge_count[5]),
	.D(N41),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[3]  (
	.SI(edge_count[2]),
	.SE(test_se),
	.RN(RST),
	.Q(edge_count[3]),
	.D(N39),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[2]  (
	.SI(edge_count[1]),
	.SE(test_se),
	.RN(RST),
	.Q(edge_count[2]),
	.D(N38),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[0]  (
	.SI(bit_count[3]),
	.SE(test_se),
	.RN(RST),
	.Q(edge_count[0]),
	.D(N36),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[4]  (
	.SI(edge_count[3]),
	.SE(test_se),
	.RN(RST),
	.Q(edge_count[4]),
	.D(N40),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[1]  (
	.SI(edge_count[0]),
	.SE(FE_OFN14_SE),
	.RN(RST),
	.Q(edge_count[1]),
	.D(N37),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_count_reg[3]  (
	.SI(bit_count[2]),
	.SE(test_se),
	.RN(RST),
	.Q(bit_count[3]),
	.D(n28),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_count_reg[2]  (
	.SI(bit_count[1]),
	.SE(test_se),
	.RN(RST),
	.Q(bit_count[2]),
	.D(n29),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_count_reg[1]  (
	.SI(bit_count[0]),
	.SE(test_se),
	.RN(RST),
	.Q(bit_count[1]),
	.D(n30),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_count_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(bit_count[0]),
	.D(n31),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U6 (
	.Y(n34),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U7 (
	.Y(n27),
	.B(N14),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U15 (
	.Y(n23),
	.C(n38),
	.B(n36),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U16 (
	.Y(n26),
	.B0(n27),
	.A1(edge_count_en),
	.A0(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n40),
	.A(edge_count_en), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U18 (
	.Y(N37),
	.B(n27),
	.A(N21), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U19 (
	.Y(N38),
	.B(n27),
	.A(N22), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U20 (
	.Y(N39),
	.B(n27),
	.A(N23), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U21 (
	.Y(N40),
	.B(n27),
	.A(N24), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U22 (
	.Y(n31),
	.B1(n34),
	.B0(n36),
	.A2(n27),
	.A1(bit_count[0]),
	.A0(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U23 (
	.Y(n29),
	.B1(n38),
	.B0(n25),
	.A2(n37),
	.A1(bit_count[2]),
	.A0(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X2M U24 (
	.Y(n25),
	.B0(n26),
	.A1(bit_count[1]),
	.A0(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U25 (
	.Y(n28),
	.B1(n40),
	.B0(n22),
	.A1(n34),
	.A0(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U26 (
	.Y(n22),
	.B1(n35),
	.B0(bit_count[3]),
	.A2(N14),
	.A1(n39),
	.A0(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U27 (
	.Y(n35),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U28 (
	.Y(n39),
	.A(bit_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U29 (
	.Y(n30),
	.B1(n24),
	.B0(bit_count[1]),
	.A1(n37),
	.A0(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U30 (
	.Y(n24),
	.C(edge_count_en),
	.B(n34),
	.A(bit_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U31 (
	.Y(n36),
	.A(bit_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U32 (
	.Y(n37),
	.A(bit_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U33 (
	.Y(n38),
	.A(bit_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U34 (
	.Y(N7),
	.A(Prescale[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U35 (
	.S(N21),
	.CO(\add_27/carry[2] ),
	.B(edge_count[0]),
	.A(edge_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U36 (
	.S(N22),
	.CO(\add_27/carry[3] ),
	.B(\add_27/carry[2] ),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U37 (
	.S(N23),
	.CO(\add_27/carry[4] ),
	.B(\add_27/carry[3] ),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U38 (
	.Y(N41),
	.B(n27),
	.A(N25), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U39 (
	.Y(N36),
	.B(n27),
	.A(N20), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U40 (
	.Y(N20),
	.A(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U41 (
	.S(N24),
	.CO(\add_27/carry[5] ),
	.B(\add_27/carry[4] ),
	.A(edge_count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U42 (
	.Y(n1),
	.B(N7),
	.AN(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U43 (
	.Y(N8),
	.B0(n1),
	.A1N(Prescale[1]),
	.A0N(Prescale[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U44 (
	.Y(n2),
	.B(Prescale[2]),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U45 (
	.Y(N9),
	.B0(n2),
	.A1N(Prescale[2]),
	.A0N(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U46 (
	.Y(n3),
	.B(Prescale[3]),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U47 (
	.Y(N10),
	.B0(n3),
	.A1N(Prescale[3]),
	.A0N(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U48 (
	.Y(n4),
	.B(Prescale[4]),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U49 (
	.Y(N11),
	.B0(n4),
	.A1N(Prescale[4]),
	.A0N(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U50 (
	.Y(N13),
	.B(Prescale[5]),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U51 (
	.Y(N12),
	.B0(N13),
	.A1(Prescale[5]),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U52 (
	.Y(N25),
	.B(edge_count[5]),
	.A(\add_27/carry[5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U53 (
	.Y(n15),
	.B(edge_count[0]),
	.AN(N7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U54 (
	.Y(n19),
	.B1(n15),
	.B0(N8),
	.A1N(edge_count[1]),
	.A0(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U55 (
	.Y(n18),
	.B(edge_count[5]),
	.A(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U56 (
	.Y(n16),
	.B(N7),
	.AN(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U57 (
	.Y(n17),
	.B1(n16),
	.B0(edge_count[1]),
	.A1N(N8),
	.A0(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U58 (
	.Y(n33),
	.D(n17),
	.C(n18),
	.B(n19),
	.AN(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U59 (
	.Y(n32),
	.B(edge_count[4]),
	.A(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U60 (
	.Y(n21),
	.B(edge_count[2]),
	.A(N9), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U61 (
	.Y(n20),
	.B(edge_count[3]),
	.A(N10), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U62 (
	.Y(N14),
	.D(n20),
	.C(n21),
	.B(n32),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Data_Sampling_test_1 (
	CLK, 
	RST, 
	Data_samp_en, 
	RX_IN, 
	Prescale, 
	edge_count, 
	Sampled_Bit, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input Data_samp_en;
   input RX_IN;
   input [5:0] Prescale;
   input [5:0] edge_count;
   output Sampled_Bit;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire sampled_bit_1;
   wire sampled_bit_2;
   wire sampled_bit_3;
   wire N7;
   wire N8;
   wire N9;
   wire N10;
   wire N11;
   wire N12;
   wire N13;
   wire N16;
   wire N17;
   wire N18;
   wire N19;
   wire N20;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire \add_33/carry[4] ;
   wire \add_33/carry[3] ;
   wire \add_33/carry[2] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;

   assign test_so = sampled_bit_3 ;

   // Module instantiations
   SDFFRQX2M sampled_bit_3_reg (
	.SI(sampled_bit_2),
	.SE(test_se),
	.RN(RST),
	.Q(sampled_bit_3),
	.D(n30),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M sampled_bit_1_reg (
	.SI(Sampled_Bit),
	.SE(test_se),
	.RN(RST),
	.Q(sampled_bit_1),
	.D(n31),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M sampled_bit_2_reg (
	.SI(sampled_bit_1),
	.SE(test_se),
	.RN(RST),
	.Q(sampled_bit_2),
	.D(n32),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M Sampled_Bit_reg (
	.SI(edge_count[5]),
	.SE(test_se),
	.RN(RST),
	.Q(Sampled_Bit),
	.D(n29),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U4 (
	.Y(n37),
	.B(Prescale[1]),
	.A(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(N7),
	.A(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U6 (
	.S(N18),
	.CO(\add_33/carry[4] ),
	.B(\add_33/carry[3] ),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U7 (
	.S(N16),
	.CO(\add_33/carry[2] ),
	.B(Prescale[1]),
	.A(Prescale[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U8 (
	.S(N17),
	.CO(\add_33/carry[3] ),
	.B(\add_33/carry[2] ),
	.A(Prescale[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U12 (
	.S(N19),
	.CO(N20),
	.B(\add_33/carry[4] ),
	.A(Prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U13 (
	.Y(n1),
	.B(N7),
	.AN(Prescale[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U14 (
	.Y(N8),
	.B0(n1),
	.A1N(Prescale[2]),
	.A0N(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U15 (
	.Y(n2),
	.B(Prescale[3]),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U16 (
	.Y(N9),
	.B0(n2),
	.A1N(Prescale[3]),
	.A0N(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U17 (
	.Y(N10),
	.B(n2),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U18 (
	.Y(N12),
	.C(n2),
	.B(Prescale[5]),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U19 (
	.Y(n3),
	.B0(Prescale[5]),
	.A1(n2),
	.A0(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U20 (
	.Y(N11),
	.B(n3),
	.AN(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U21 (
	.Y(n4),
	.B(N7),
	.AN(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U22 (
	.Y(n7),
	.B1(n4),
	.B0(edge_count[1]),
	.A1N(N8),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U23 (
	.Y(n5),
	.B(edge_count[0]),
	.AN(N7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U24 (
	.Y(n6),
	.B1(n5),
	.B0(N8),
	.A1N(edge_count[1]),
	.A0(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BBX1M U25 (
	.Y(n15),
	.D(n6),
	.C(n7),
	.BN(edge_count[5]),
	.AN(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U26 (
	.Y(n10),
	.B(edge_count[4]),
	.A(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U27 (
	.Y(n9),
	.B(edge_count[2]),
	.A(N9), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U28 (
	.Y(n8),
	.B(edge_count[3]),
	.A(N10), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U29 (
	.Y(N13),
	.D(n8),
	.C(n9),
	.B(n10),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U30 (
	.Y(n32),
	.S0(n18),
	.B(n17),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U31 (
	.Y(n16),
	.B(Data_samp_en),
	.A(sampled_bit_2), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U32 (
	.Y(n31),
	.S0(n20),
	.B(n19),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U33 (
	.Y(n19),
	.B(Data_samp_en),
	.A(sampled_bit_1), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U34 (
	.Y(n30),
	.S0(n22),
	.B(n21),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X1M U35 (
	.Y(n22),
	.B0(n25),
	.A2(n24),
	.A1(n20),
	.A0(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U36 (
	.Y(n20),
	.A(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U37 (
	.Y(n21),
	.A(sampled_bit_3), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U38 (
	.Y(n17),
	.B(Data_samp_en),
	.A(RX_IN), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U39 (
	.Y(n29),
	.B(n26),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U40 (
	.Y(n26),
	.S0(n28),
	.B(n27),
	.A(Sampled_Bit), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U41 (
	.Y(n28),
	.C(n24),
	.B(N13),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X1M U42 (
	.Y(n24),
	.D(n36),
	.C(n35),
	.B(n34),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U43 (
	.Y(n36),
	.C(n39),
	.B(n38),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U44 (
	.Y(n39),
	.B(N19),
	.A(edge_count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U45 (
	.Y(n38),
	.B(N16),
	.A(edge_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U46 (
	.Y(n35),
	.B(N17),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U47 (
	.Y(n34),
	.B(N18),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U48 (
	.Y(n33),
	.B(N20),
	.A(edge_count[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U49 (
	.Y(n18),
	.B(N13),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U50 (
	.Y(n23),
	.D(n43),
	.C(n42),
	.B(n41),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U51 (
	.Y(n43),
	.C(n45),
	.B(edge_count[5]),
	.A(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U52 (
	.Y(n45),
	.B(Prescale[1]),
	.A(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U53 (
	.Y(n44),
	.B(Prescale[5]),
	.A(edge_count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U54 (
	.Y(n42),
	.B(Prescale[3]),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U55 (
	.Y(n41),
	.B(Prescale[4]),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U56 (
	.Y(n40),
	.B(Prescale[2]),
	.A(edge_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U57 (
	.Y(n27),
	.B0(n46),
	.A1N(sampled_bit_1),
	.A0N(sampled_bit_2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U58 (
	.Y(n46),
	.B0(sampled_bit_3),
	.A1(sampled_bit_2),
	.A0(sampled_bit_1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U59 (
	.Y(n25),
	.A(Data_samp_en), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Start_Check_test_1 (
	CLK, 
	RST, 
	start_en, 
	Sampled_Bit, 
	Start_glitch, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input start_en;
   input Sampled_Bit;
   output Start_glitch;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N4;

   // Module instantiations
   SDFFRQX2M Start_glitch_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(Start_glitch),
	.D(N4),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U4 (
	.Y(N4),
	.B(Sampled_Bit),
	.A(start_en), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Stop_Check_test_1 (
	CLK, 
	RST, 
	stop_en, 
	Sampled_Bit, 
	Stop_error, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input stop_en;
   input Sampled_Bit;
   output Stop_error;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n3;

   // Module instantiations
   SDFFRQX4M Stop_error_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(Stop_error),
	.D(n3),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U2 (
	.Y(n3),
	.B1(stop_en),
	.B0(Sampled_Bit),
	.A1N(stop_en),
	.A0N(Stop_error), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Deserializer_test_1 (
	CLK, 
	RST, 
	desrializer_en, 
	Sampled_Bit, 
	DATA_VALID, 
	bit_count, 
	parity_flag, 
	P_DATA, 
	test_si, 
	test_se, 
	FE_OFN11_SE, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input desrializer_en;
   input Sampled_Bit;
   input DATA_VALID;
   input [3:0] bit_count;
   output parity_flag;
   output [7:0] P_DATA;
   input test_si;
   input test_se;
   input FE_OFN11_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire [7:0] DATA;

   // Module instantiations
   SDFFQX2M \DATA_reg[5]  (
	.SI(DATA[4]),
	.SE(FE_OFN11_SE),
	.Q(DATA[5]),
	.D(n41),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \DATA_reg[1]  (
	.SI(DATA[0]),
	.SE(test_se),
	.Q(DATA[1]),
	.D(n37),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \DATA_reg[4]  (
	.SI(DATA[3]),
	.SE(test_se),
	.Q(DATA[4]),
	.D(n40),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \DATA_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.Q(DATA[0]),
	.D(n36),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M parity_flag_reg (
	.SI(DATA[7]),
	.SE(FE_OFN11_SE),
	.RN(RST),
	.Q(parity_flag),
	.D(n35),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \DATA_reg[2]  (
	.SI(DATA[1]),
	.SE(test_se),
	.Q(DATA[2]),
	.D(n38),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \DATA_reg[3]  (
	.SI(DATA[2]),
	.SE(test_se),
	.Q(DATA[3]),
	.D(n39),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \DATA_reg[6]  (
	.SI(DATA[5]),
	.SE(FE_OFN11_SE),
	.Q(DATA[6]),
	.D(n42),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \DATA_reg[7]  (
	.SI(DATA[6]),
	.SE(FE_OFN11_SE),
	.Q(DATA[7]),
	.D(n43),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(n10),
	.A(RST), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U13 (
	.Y(n32),
	.B(DATA_VALID),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U14 (
	.Y(n11),
	.A(DATA_VALID), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U15 (
	.Y(n28),
	.B(n16),
	.AN(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U16 (
	.Y(n12),
	.A(desrializer_en), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3BX2M U17 (
	.Y(n25),
	.C(n15),
	.B(bit_count[2]),
	.AN(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3BX2M U18 (
	.Y(n23),
	.C(bit_count[3]),
	.B(n10),
	.AN(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U19 (
	.Y(n21),
	.B(DATA[3]),
	.A(DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n14),
	.A(bit_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n15),
	.A(bit_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n13),
	.A(Sampled_Bit), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U23 (
	.Y(n35),
	.B1(n12),
	.B0(n17),
	.A1N(n12),
	.A0N(parity_flag), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U24 (
	.Y(n17),
	.B(n19),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U25 (
	.Y(n19),
	.C(n20),
	.B(DATA[4]),
	.A(DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U26 (
	.Y(n18),
	.C(n21),
	.B(DATA[0]),
	.A(DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U27 (
	.Y(n39),
	.B1(n27),
	.B0(n13),
	.A1N(DATA[3]),
	.A0N(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U28 (
	.Y(n27),
	.C(n28),
	.B(n15),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U29 (
	.Y(n37),
	.B1(n24),
	.B0(n13),
	.A1N(DATA[1]),
	.A0N(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U30 (
	.Y(n24),
	.B(n14),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U31 (
	.Y(n38),
	.B1(n26),
	.B0(n13),
	.A1N(DATA[2]),
	.A0N(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U32 (
	.Y(n26),
	.B(bit_count[0]),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U33 (
	.Y(n36),
	.B1(n13),
	.B0(n22),
	.A1N(DATA[0]),
	.A0N(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U34 (
	.Y(n22),
	.D(n16),
	.C(n15),
	.B(n23),
	.A(bit_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U35 (
	.Y(n40),
	.B1(n29),
	.B0(n13),
	.A1N(DATA[4]),
	.A0N(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U36 (
	.Y(n29),
	.C(n28),
	.B(n15),
	.A(bit_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U37 (
	.Y(n41),
	.B1(n30),
	.B0(n13),
	.A1N(DATA[5]),
	.A0N(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U38 (
	.Y(n30),
	.C(n28),
	.B(n14),
	.A(bit_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U39 (
	.Y(n42),
	.B1(n31),
	.B0(n13),
	.A1N(DATA[6]),
	.A0N(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U40 (
	.Y(n31),
	.C(n28),
	.B(bit_count[0]),
	.A(bit_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U41 (
	.Y(n43),
	.B1(n33),
	.B0(n13),
	.A1N(DATA[7]),
	.A0N(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U42 (
	.Y(n33),
	.D(n34),
	.C(bit_count[3]),
	.B(RST),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U43 (
	.Y(n34),
	.C(bit_count[1]),
	.B(bit_count[2]),
	.A(bit_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U44 (
	.Y(n16),
	.A(bit_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U45 (
	.Y(P_DATA[0]),
	.B(DATA_VALID),
	.A(DATA[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U46 (
	.Y(P_DATA[1]),
	.B(DATA_VALID),
	.A(DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U47 (
	.Y(P_DATA[2]),
	.B(n11),
	.AN(DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U48 (
	.Y(P_DATA[3]),
	.B(n11),
	.AN(DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U49 (
	.Y(P_DATA[4]),
	.B(DATA_VALID),
	.A(DATA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U50 (
	.Y(P_DATA[5]),
	.B(DATA_VALID),
	.A(DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U51 (
	.Y(P_DATA[6]),
	.B(n11),
	.AN(DATA[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U52 (
	.Y(P_DATA[7]),
	.B(DATA_VALID),
	.A(DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U53 (
	.Y(n20),
	.B(DATA[6]),
	.A(DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Parity_Check_test_1 (
	CLK, 
	RST, 
	Parity_type, 
	parity_check_en, 
	Sampled_Bit, 
	parity_flag, 
	Parity_error, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input Parity_type;
   input parity_check_en;
   input Sampled_Bit;
   input parity_flag;
   output Parity_error;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n3;

   // Module instantiations
   SDFFRQX4M Parity_error_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(Parity_error),
	.D(n3),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U3 (
	.Y(n3),
	.B1(n1),
	.B0(parity_check_en),
	.A1N(parity_check_en),
	.A0(Parity_error), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U4 (
	.Y(n1),
	.C(Parity_type),
	.B(Sampled_Bit),
	.A(parity_flag), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_TX_TOP_DATA_WIDTH8_test_1 (
	CLK, 
	RST, 
	party_en, 
	data_valid, 
	party_typ, 
	P_DATA, 
	busy, 
	Tx_OUT, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN13_SE, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input party_en;
   input data_valid;
   input party_typ;
   input [7:0] P_DATA;
   output busy;
   output Tx_OUT;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN13_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire ser_done;
   wire ser_en;
   wire ser_data;
   wire party_bit;
   wire n2;
   wire [2:0] mux_sel;

   // Module instantiations
   serializer_DATA_WIDTH8_test_1 serial (
	.P_DATA({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }),
	.ser_en(ser_en),
	.RST(RST),
	.CLK(CLK),
	.data_valid(data_valid),
	.ser_done(ser_done),
	.ser_data(ser_data),
	.test_si(n2),
	.test_so(test_so),
	.test_se(test_se),
	.FE_OFN13_SE(FE_OFN13_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   FSM_TX_test_1 FSM (
	.CLK(CLK),
	.RST(RST),
	.party_en(party_en),
	.ser_done(ser_done),
	.data_valid(data_valid),
	.busy(busy),
	.ser_en(ser_en),
	.mux_sel({ mux_sel[2],
		mux_sel[1],
		mux_sel[0] }),
	.test_si(test_si),
	.test_so(n2),
	.test_se(test_se),
	.FE_OFN13_SE(FE_OFN13_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   parity_calc_DATA_WIDTH8 parity (
	.party_typ(party_typ),
	.data_valid(data_valid),
	.CLK(1'b0),
	.RST(1'b0),
	.busy(1'b0),
	.P_DATA({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }),
	.party_bit(party_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   MUX MUX (
	.mux_sel({ mux_sel[2],
		mux_sel[1],
		mux_sel[0] }),
	.ser_data(ser_data),
	.party_bit(party_bit),
	.Tx_OUT(Tx_OUT), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module serializer_DATA_WIDTH8_test_1 (
	P_DATA, 
	ser_en, 
	RST, 
	CLK, 
	data_valid, 
	ser_done, 
	ser_data, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN13_SE, 
	VDD, 
	VSS);
   input [7:0] P_DATA;
   input ser_en;
   input RST;
   input CLK;
   input data_valid;
   output ser_done;
   output ser_data;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN13_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N3;
   wire N4;
   wire N5;
   wire N16;
   wire N17;
   wire N18;
   wire N24;
   wire n2;
   wire n7;
   wire n8;
   wire n10;
   wire n12;
   wire n14;
   wire n16;
   wire n18;
   wire n20;
   wire n22;
   wire n24;
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n28;
   wire n29;
   wire [7:0] P_DATA_COMP;

   assign test_so = N5 ;

   // Module instantiations
   SDFFRQX2M \P_DATA_COMP_reg[5]  (
	.SI(P_DATA_COMP[4]),
	.SE(FE_OFN13_SE),
	.RN(RST),
	.Q(P_DATA_COMP[5]),
	.D(n20),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_COMP_reg[1]  (
	.SI(P_DATA_COMP[0]),
	.SE(FE_OFN13_SE),
	.RN(RST),
	.Q(P_DATA_COMP[1]),
	.D(n12),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_COMP_reg[7]  (
	.SI(P_DATA_COMP[6]),
	.SE(FE_OFN13_SE),
	.RN(RST),
	.Q(P_DATA_COMP[7]),
	.D(n24),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_COMP_reg[3]  (
	.SI(P_DATA_COMP[2]),
	.SE(FE_OFN13_SE),
	.RN(RST),
	.Q(P_DATA_COMP[3]),
	.D(n16),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_COMP_reg[6]  (
	.SI(P_DATA_COMP[5]),
	.SE(FE_OFN13_SE),
	.RN(RST),
	.Q(P_DATA_COMP[6]),
	.D(n22),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_COMP_reg[2]  (
	.SI(P_DATA_COMP[1]),
	.SE(FE_OFN13_SE),
	.RN(RST),
	.Q(P_DATA_COMP[2]),
	.D(n14),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_COMP_reg[4]  (
	.SI(P_DATA_COMP[3]),
	.SE(FE_OFN13_SE),
	.RN(RST),
	.Q(P_DATA_COMP[4]),
	.D(n18),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_COMP_reg[0]  (
	.SI(test_si),
	.SE(FE_OFN13_SE),
	.RN(RST),
	.Q(P_DATA_COMP[0]),
	.D(n10),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[1]  (
	.SI(N3),
	.SE(FE_OFN13_SE),
	.RN(RST),
	.Q(N4),
	.D(N17),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[2]  (
	.SI(N4),
	.SE(test_se),
	.RN(RST),
	.Q(N5),
	.D(N18),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[0]  (
	.SI(P_DATA_COMP[7]),
	.SE(FE_OFN13_SE),
	.RN(RST),
	.Q(N3),
	.D(N16),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(n5),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U4 (
	.Y(n2),
	.D(n29),
	.C(n28),
	.B(n6),
	.A(data_valid), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U5 (
	.Y(N17),
	.C0(n7),
	.B0(n4),
	.A1(n28),
	.A0(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U6 (
	.Y(n7),
	.B(n6),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U7 (
	.Y(n4),
	.A(ser_en), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U8 (
	.Y(ser_data),
	.B(n4),
	.AN(N24), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U9 (
	.Y(N24),
	.S0(N5),
	.B(n1),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U10 (
	.Y(n1),
	.S1(N4),
	.S0(N3),
	.D(P_DATA_COMP[7]),
	.C(P_DATA_COMP[6]),
	.B(P_DATA_COMP[5]),
	.A(P_DATA_COMP[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U11 (
	.Y(n3),
	.S1(N4),
	.S0(N3),
	.D(P_DATA_COMP[3]),
	.C(P_DATA_COMP[2]),
	.B(P_DATA_COMP[1]),
	.A(P_DATA_COMP[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U12 (
	.Y(N18),
	.B1(n4),
	.B0(n8),
	.A1N(N16),
	.A0N(N5), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U13 (
	.Y(n8),
	.B1(n28),
	.B0(N5),
	.A1(n29),
	.A0(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U14 (
	.Y(N16),
	.B(N3),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U15 (
	.Y(n6),
	.A(N3), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U16 (
	.Y(n28),
	.A(N4), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n29),
	.A(N5), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U18 (
	.Y(ser_done),
	.B(N5),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U19 (
	.Y(n10),
	.B1(n5),
	.B0(P_DATA[0]),
	.A1(n2),
	.A0(P_DATA_COMP[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U20 (
	.Y(n12),
	.B1(n5),
	.B0(P_DATA[1]),
	.A1(n2),
	.A0(P_DATA_COMP[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U21 (
	.Y(n14),
	.B1(n5),
	.B0(P_DATA[2]),
	.A1(n2),
	.A0(P_DATA_COMP[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U22 (
	.Y(n16),
	.B1(n5),
	.B0(P_DATA[3]),
	.A1(n2),
	.A0(P_DATA_COMP[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U23 (
	.Y(n18),
	.B1(n5),
	.B0(P_DATA[4]),
	.A1(n2),
	.A0(P_DATA_COMP[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U35 (
	.Y(n20),
	.B1(n5),
	.B0(P_DATA[5]),
	.A1(n2),
	.A0(P_DATA_COMP[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U36 (
	.Y(n22),
	.B1(n5),
	.B0(P_DATA[6]),
	.A1(n2),
	.A0(P_DATA_COMP[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U37 (
	.Y(n24),
	.B1(n5),
	.B0(P_DATA[7]),
	.A1(n2),
	.A0(P_DATA_COMP[7]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FSM_TX_test_1 (
	CLK, 
	RST, 
	party_en, 
	ser_done, 
	data_valid, 
	busy, 
	ser_en, 
	mux_sel, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN13_SE, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input party_en;
   input ser_done;
   input data_valid;
   output busy;
   output ser_en;
   output [2:0] mux_sel;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN13_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n5;
   wire n6;
   wire [2:0] current_state;
   wire [2:0] next_state;

   assign test_so = current_state[2] ;

   // Module instantiations
   SDFFRQX2M \current_state_reg[1]  (
	.SI(current_state[0]),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[1]),
	.D(next_state[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[0]  (
	.SI(test_si),
	.SE(FE_OFN13_SE),
	.RN(RST),
	.Q(current_state[0]),
	.D(next_state[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[2]  (
	.SI(current_state[1]),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[2]),
	.D(next_state[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U6 (
	.Y(mux_sel[2]),
	.A(busy), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U7 (
	.Y(busy),
	.B1(n5),
	.B0(n6),
	.A1(current_state[2]),
	.A0(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U8 (
	.Y(ser_en),
	.C(n6),
	.B(current_state[2]),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U9 (
	.Y(n8),
	.B0(mux_sel[1]),
	.A1(current_state[0]),
	.A0(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U10 (
	.Y(mux_sel[1]),
	.B(current_state[0]),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21BX1M U11 (
	.Y(next_state[1]),
	.B0N(ser_en),
	.A1(n8),
	.A0(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X1M U12 (
	.Y(next_state[2]),
	.B0(current_state[2]),
	.A1N(mux_sel[1]),
	.A0(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U13 (
	.Y(n7),
	.C(ser_done),
	.B(current_state[1]),
	.AN(party_en), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U14 (
	.Y(next_state[0]),
	.B0(current_state[2]),
	.A1(n10),
	.A0(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U15 (
	.Y(n9),
	.B(n5),
	.A(ser_done), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U16 (
	.Y(n10),
	.B0(n6),
	.A1(data_valid),
	.A0(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n6),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(n5),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U19 (
	.Y(mux_sel[0]),
	.B(current_state[2]),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module parity_calc_DATA_WIDTH8 (
	party_typ, 
	data_valid, 
	CLK, 
	RST, 
	busy, 
	P_DATA, 
	party_bit, 
	VDD, 
	VSS);
   input party_typ;
   input data_valid;
   input CLK;
   input RST;
   input busy;
   input [7:0] P_DATA;
   output party_bit;
   inout VDD;
   inout VSS;

   // Internal wires
   wire LTIE_LTIELO_NET;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n8;

   // Module instantiations
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M party_bit_reg (
	.SI(LTIE_LTIELO_NET),
	.SE(LTIE_LTIELO_NET),
	.RN(LTIE_LTIELO_NET),
	.Q(party_bit),
	.D(n8),
	.CK(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U2 (
	.Y(n4),
	.C(n5),
	.B(P_DATA[0]),
	.A(P_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U3 (
	.Y(n5),
	.B(P_DATA[2]),
	.A(P_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U4 (
	.Y(n8),
	.B1(n2),
	.B0(n1),
	.A1N(n2),
	.A0N(party_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U5 (
	.Y(n2),
	.B(data_valid),
	.AN(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U6 (
	.Y(n1),
	.C(n4),
	.B(party_typ),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U7 (
	.Y(n3),
	.C(n6),
	.B(P_DATA[4]),
	.A(P_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U8 (
	.Y(n6),
	.B(P_DATA[6]),
	.A(P_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module MUX (
	mux_sel, 
	ser_data, 
	party_bit, 
	Tx_OUT, 
	VDD, 
	VSS);
   input [2:0] mux_sel;
   input ser_data;
   input party_bit;
   output Tx_OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n2;

   // Module instantiations
   NAND3BX4M U3 (
	.Y(Tx_OUT),
	.C(n2),
	.B(n1),
	.AN(mux_sel[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U4 (
	.Y(n2),
	.B(mux_sel[0]),
	.A(ser_data), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U5 (
	.Y(n1),
	.B0(mux_sel[1]),
	.A1(party_bit),
	.A0(mux_sel[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SYSTEM_CONTROL_DATA_WIDTH8_test_1 (
	REF_CLK, 
	RST_SYNC_2, 
	pulse_gen, 
	W_FULL, 
	R_DATA_VALID, 
	ALU_OUT_VALID, 
	SYNC_BUS, 
	R_REG_DATA, 
	ALU_OUT, 
	WINC, 
	W_REG_EN, 
	R_REG_EN, 
	ALU_EN, 
	CLK_GATE_EN, 
	div_en, 
	W_DATA, 
	W_REG_DATA, 
	REG_ADDRESS, 
	ALU_FUNC, 
	test_si, 
	test_so, 
	test_se, 
	scanclkref__L7_N1, 
	VDD, 
	VSS);
   input REF_CLK;
   input RST_SYNC_2;
   input pulse_gen;
   input W_FULL;
   input R_DATA_VALID;
   input ALU_OUT_VALID;
   input [7:0] SYNC_BUS;
   input [7:0] R_REG_DATA;
   input [15:0] ALU_OUT;
   output WINC;
   output W_REG_EN;
   output R_REG_EN;
   output ALU_EN;
   output CLK_GATE_EN;
   output div_en;
   output [7:0] W_DATA;
   output [7:0] W_REG_DATA;
   output [3:0] REG_ADDRESS;
   output [3:0] ALU_FUNC;
   input test_si;
   output test_so;
   input test_se;
   input scanclkref__L7_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN9_REG_ADDRESS_1_;
   wire FE_OFN8_REG_ADDRESS_3_;
   wire FE_OFN7_REG_ADDRESS_2_;
   wire \comb_reg_address[0] ;
   wire n27;
   wire n28;
   wire n29;
   wire n41;
   wire n42;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n69;
   wire n70;
   wire n71;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n16;
   wire n17;
   wire n18;
   wire n22;
   wire n23;
   wire n24;
   wire n26;
   wire n30;
   wire n32;
   wire n33;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n43;
   wire n68;
   wire n72;
   wire n81;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire [3:0] current_state;
   wire [2:0] next_state;
   wire [7:0] W_DATA_2;

   assign div_en = 1'b1 ;
   assign test_so = current_state[2] ;

   // Module instantiations
   BUFX2M FE_OFC9_REG_ADDRESS_1_ (
	.Y(REG_ADDRESS[1]),
	.A(FE_OFN9_REG_ADDRESS_1_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M FE_OFC8_REG_ADDRESS_3_ (
	.Y(REG_ADDRESS[3]),
	.A(FE_OFN8_REG_ADDRESS_3_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M FE_OFC7_REG_ADDRESS_2_ (
	.Y(REG_ADDRESS[2]),
	.A(FE_OFN7_REG_ADDRESS_2_), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \comb_reg_address_reg[3]  (
	.SI(n102),
	.SE(test_se),
	.RN(RST_SYNC_2),
	.QN(n27),
	.Q(n101),
	.D(n90),
	.CK(scanclkref__L7_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \comb_reg_address_reg[2]  (
	.SI(n103),
	.SE(test_se),
	.RN(RST_SYNC_2),
	.QN(n28),
	.Q(n102),
	.D(n89),
	.CK(scanclkref__L7_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \comb_reg_address_reg[1]  (
	.SI(\comb_reg_address[0] ),
	.SE(test_se),
	.RN(RST_SYNC_2),
	.QN(n29),
	.Q(n103),
	.D(n88),
	.CK(scanclkref__L7_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \W_DATA_2_reg[7]  (
	.SI(W_DATA_2[6]),
	.SE(test_se),
	.RN(RST_SYNC_2),
	.Q(W_DATA_2[7]),
	.D(n98),
	.CK(REF_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \W_DATA_2_reg[6]  (
	.SI(W_DATA_2[5]),
	.SE(test_se),
	.RN(RST_SYNC_2),
	.Q(W_DATA_2[6]),
	.D(n97),
	.CK(REF_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \W_DATA_2_reg[5]  (
	.SI(W_DATA_2[4]),
	.SE(test_se),
	.RN(RST_SYNC_2),
	.Q(W_DATA_2[5]),
	.D(n96),
	.CK(REF_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \W_DATA_2_reg[4]  (
	.SI(W_DATA_2[3]),
	.SE(test_se),
	.RN(RST_SYNC_2),
	.Q(W_DATA_2[4]),
	.D(n95),
	.CK(REF_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \W_DATA_2_reg[3]  (
	.SI(W_DATA_2[2]),
	.SE(test_se),
	.RN(RST_SYNC_2),
	.Q(W_DATA_2[3]),
	.D(n94),
	.CK(REF_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \W_DATA_2_reg[2]  (
	.SI(W_DATA_2[1]),
	.SE(test_se),
	.RN(RST_SYNC_2),
	.Q(W_DATA_2[2]),
	.D(n93),
	.CK(REF_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \W_DATA_2_reg[1]  (
	.SI(W_DATA_2[0]),
	.SE(test_se),
	.RN(RST_SYNC_2),
	.Q(W_DATA_2[1]),
	.D(n92),
	.CK(REF_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \W_DATA_2_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST_SYNC_2),
	.Q(W_DATA_2[0]),
	.D(n91),
	.CK(REF_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \comb_reg_address_reg[0]  (
	.SI(W_DATA_2[7]),
	.SE(test_se),
	.RN(RST_SYNC_2),
	.Q(\comb_reg_address[0] ),
	.D(n87),
	.CK(scanclkref__L7_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[1]  (
	.SI(current_state[0]),
	.SE(test_se),
	.RN(RST_SYNC_2),
	.Q(current_state[1]),
	.D(next_state[1]),
	.CK(REF_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[2]  (
	.SI(current_state[1]),
	.SE(test_se),
	.RN(RST_SYNC_2),
	.Q(current_state[2]),
	.D(next_state[2]),
	.CK(REF_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[0]  (
	.SI(n101),
	.SE(test_se),
	.RN(RST_SYNC_2),
	.Q(current_state[0]),
	.D(next_state[0]),
	.CK(scanclkref__L7_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U18 (
	.Y(ALU_FUNC[2]),
	.B(n86),
	.A(n81), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U19 (
	.Y(ALU_FUNC[0]),
	.B(n86),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U20 (
	.Y(FE_OFN7_REG_ADDRESS_2_),
	.B1(n84),
	.B0(n28),
	.A1(n83),
	.A0(n81), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n24),
	.A(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U23 (
	.Y(CLK_GATE_EN),
	.B(n30),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U24 (
	.Y(n30),
	.A(n71), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U25 (
	.Y(n23),
	.A(W_FULL), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U26 (
	.Y(n67),
	.C(n38),
	.B(n32),
	.A(n60), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U27 (
	.Y(n45),
	.D(n60),
	.C(n72),
	.B(n39),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U28 (
	.Y(W_REG_DATA[0]),
	.B(n70),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U29 (
	.Y(W_REG_DATA[2]),
	.B(n70),
	.A(n81), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U30 (
	.Y(W_REG_DATA[3]),
	.B(n70),
	.A(n72), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U31 (
	.Y(W_REG_DATA[4]),
	.B(n70),
	.A(n68), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U32 (
	.Y(W_REG_DATA[5]),
	.B(n70),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U33 (
	.Y(W_REG_DATA[6]),
	.B(n70),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U34 (
	.Y(W_REG_DATA[7]),
	.B(n70),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U35 (
	.Y(W_REG_DATA[1]),
	.B(n70),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U36 (
	.Y(ALU_FUNC[1]),
	.B(n86),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21BX1M U37 (
	.Y(n51),
	.B0N(n61),
	.A1(n60),
	.A0(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U38 (
	.Y(WINC),
	.B0(n82),
	.A1(n33),
	.A0(n62), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U39 (
	.Y(n82),
	.B0(n23),
	.A1(n16),
	.A0(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4BX1M U40 (
	.Y(n58),
	.D(n99),
	.C(n43),
	.B(n59),
	.AN(n45), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U41 (
	.Y(n59),
	.D(n32),
	.C(n40),
	.B(n81),
	.A(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U42 (
	.Y(n33),
	.A(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U43 (
	.Y(n60),
	.B(n36),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U44 (
	.Y(ALU_EN),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U45 (
	.Y(ALU_FUNC[3]),
	.B(n86),
	.A(n72), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U46 (
	.Y(n35),
	.A(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U47 (
	.Y(n71),
	.B(n61),
	.A(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U48 (
	.Y(R_REG_EN),
	.A(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U49 (
	.Y(W_REG_EN),
	.A(n70), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X2M U52 (
	.Y(FE_OFN8_REG_ADDRESS_3_),
	.B1(n84),
	.B0(n27),
	.A1(n83),
	.A0(n72), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U53 (
	.Y(n49),
	.C(n37),
	.B(current_state[2]),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U54 (
	.Y(n53),
	.C(n37),
	.B(current_state[0]),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U55 (
	.Y(n64),
	.C(n37),
	.B(current_state[2]),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U56 (
	.Y(n50),
	.B1(n23),
	.B0(n66),
	.A1N(n64),
	.A0(n65), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U57 (
	.Y(n65),
	.B(W_FULL),
	.AN(R_DATA_VALID), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U58 (
	.Y(n61),
	.C(n36),
	.B(current_state[1]),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U59 (
	.Y(n63),
	.C(n36),
	.B(current_state[1]),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U60 (
	.Y(next_state[2]),
	.C0(n26),
	.B1(n23),
	.B0(n66),
	.A1(n42),
	.A0(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U61 (
	.Y(n26),
	.A(CLK_GATE_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U62 (
	.Y(n41),
	.C(n99),
	.B(n32),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U63 (
	.Y(n42),
	.D(n45),
	.C(n44),
	.B(SYNC_BUS[2]),
	.A(SYNC_BUS[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U64 (
	.Y(n86),
	.B(n53),
	.A(pulse_gen), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U65 (
	.Y(n88),
	.B1(n29),
	.B0(n67),
	.A1(n24),
	.A0(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U66 (
	.Y(n89),
	.B1(n28),
	.B0(n67),
	.A1(n24),
	.A0(n81), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U67 (
	.Y(n90),
	.B1(n27),
	.B0(n67),
	.A1(n24),
	.A0(n72), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U68 (
	.Y(n83),
	.B(n64),
	.A(pulse_gen), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U69 (
	.Y(n18),
	.B(n33),
	.AN(ALU_OUT_VALID), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U70 (
	.Y(n69),
	.B(n33),
	.AN(ALU_OUT_VALID), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U71 (
	.Y(n17),
	.B(n33),
	.AN(ALU_OUT_VALID), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U72 (
	.Y(n32),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U73 (
	.Y(n38),
	.A(pulse_gen), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U74 (
	.Y(n84),
	.B(n49),
	.A(pulse_gen), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U75 (
	.Y(n99),
	.A(SYNC_BUS[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U76 (
	.Y(n81),
	.A(SYNC_BUS[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U77 (
	.Y(n66),
	.C(current_state[1]),
	.B(current_state[0]),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U78 (
	.Y(W_DATA[0]),
	.B0(n80),
	.A1N(n16),
	.A0N(R_REG_DATA[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U79 (
	.Y(n80),
	.B1(n18),
	.B0(ALU_OUT[0]),
	.A1(n35),
	.A0(W_DATA_2[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U80 (
	.Y(W_DATA[1]),
	.B0(n79),
	.A1N(n16),
	.A0N(R_REG_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U81 (
	.Y(n79),
	.B1(n69),
	.B0(ALU_OUT[1]),
	.A1(n35),
	.A0(W_DATA_2[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U82 (
	.Y(W_DATA[2]),
	.B0(n78),
	.A1N(n16),
	.A0N(R_REG_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U83 (
	.Y(n78),
	.B1(n17),
	.B0(ALU_OUT[2]),
	.A1(n35),
	.A0(W_DATA_2[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U84 (
	.Y(W_DATA[3]),
	.B0(n77),
	.A1N(n16),
	.A0N(R_REG_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U85 (
	.Y(n77),
	.B1(n18),
	.B0(ALU_OUT[3]),
	.A1(n35),
	.A0(W_DATA_2[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U86 (
	.Y(W_DATA[4]),
	.B0(n76),
	.A1N(n16),
	.A0N(R_REG_DATA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U87 (
	.Y(n76),
	.B1(n69),
	.B0(ALU_OUT[4]),
	.A1(n35),
	.A0(W_DATA_2[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U88 (
	.Y(W_DATA[5]),
	.B0(n75),
	.A1N(n16),
	.A0N(R_REG_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U89 (
	.Y(n75),
	.B1(n17),
	.B0(ALU_OUT[5]),
	.A1(n35),
	.A0(W_DATA_2[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U90 (
	.Y(W_DATA[6]),
	.B0(n74),
	.A1N(n16),
	.A0N(R_REG_DATA[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U91 (
	.Y(n74),
	.B1(n18),
	.B0(ALU_OUT[6]),
	.A1(n35),
	.A0(W_DATA_2[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U92 (
	.Y(W_DATA[7]),
	.B0(n73),
	.A1N(n16),
	.A0N(R_REG_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U93 (
	.Y(n73),
	.B1(n69),
	.B0(ALU_OUT[7]),
	.A1(n35),
	.A0(W_DATA_2[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U94 (
	.Y(n72),
	.A(SYNC_BUS[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U95 (
	.Y(n87),
	.B1(n24),
	.B0(n100),
	.A1N(\comb_reg_address[0] ),
	.A0N(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U96 (
	.Y(n37),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U97 (
	.Y(n36),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U98 (
	.Y(n70),
	.B0(pulse_gen),
	.A1(n71),
	.A0(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U99 (
	.Y(n52),
	.B0(n68),
	.A1(n55),
	.A0(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U100 (
	.Y(n54),
	.D(n40),
	.C(n81),
	.B(SYNC_BUS[1]),
	.A(SYNC_BUS[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U101 (
	.Y(n55),
	.D(n43),
	.C(n99),
	.B(SYNC_BUS[2]),
	.A(SYNC_BUS[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U102 (
	.Y(next_state[0]),
	.B(n57),
	.A(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U103 (
	.Y(n56),
	.B0(n50),
	.A1(pulse_gen),
	.A0(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U104 (
	.Y(n57),
	.C0(n58),
	.B1(n38),
	.B0(n51),
	.A1(n53),
	.A0(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U105 (
	.Y(n22),
	.A(n62), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U106 (
	.Y(n62),
	.B(n23),
	.A(ALU_OUT_VALID), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U107 (
	.Y(n40),
	.A(SYNC_BUS[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U108 (
	.Y(n43),
	.A(SYNC_BUS[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U109 (
	.Y(n100),
	.A(SYNC_BUS[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U110 (
	.Y(n44),
	.B(SYNC_BUS[0]),
	.A(n68), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U111 (
	.Y(next_state[1]),
	.C(n46),
	.B(n48),
	.A(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U112 (
	.Y(n47),
	.B(n51),
	.A(pulse_gen), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U113 (
	.Y(n48),
	.B0(n50),
	.A1(n38),
	.A0(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U114 (
	.Y(n46),
	.B0(n53),
	.A2(n52),
	.A1(SYNC_BUS[0]),
	.A0(n45), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U115 (
	.Y(n39),
	.A(SYNC_BUS[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U116 (
	.Y(n68),
	.A(SYNC_BUS[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U117 (
	.Y(n91),
	.B1(n17),
	.B0(ALU_OUT[8]),
	.A1N(n18),
	.A0(W_DATA_2[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U118 (
	.Y(n92),
	.B1(n69),
	.B0(ALU_OUT[9]),
	.A1N(n17),
	.A0(W_DATA_2[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U119 (
	.Y(n93),
	.B1(n18),
	.B0(ALU_OUT[10]),
	.A1N(n69),
	.A0(W_DATA_2[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U120 (
	.Y(n94),
	.B1(n17),
	.B0(ALU_OUT[11]),
	.A1N(n18),
	.A0(W_DATA_2[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U121 (
	.Y(n95),
	.B1(n69),
	.B0(ALU_OUT[12]),
	.A1N(n17),
	.A0(W_DATA_2[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U122 (
	.Y(n96),
	.B1(n18),
	.B0(ALU_OUT[13]),
	.A1N(n17),
	.A0(W_DATA_2[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U123 (
	.Y(n97),
	.B1(n17),
	.B0(ALU_OUT[14]),
	.A1N(n18),
	.A0(W_DATA_2[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U124 (
	.Y(n98),
	.B1(n69),
	.B0(ALU_OUT[15]),
	.A1N(n17),
	.A0(W_DATA_2[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U125 (
	.Y(n16),
	.B(n64),
	.A(R_DATA_VALID), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U126 (
	.Y(REG_ADDRESS[0]),
	.B1(n38),
	.B0(n85),
	.A1(n83),
	.A0(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U127 (
	.Y(n85),
	.B0(n61),
	.A1(n49),
	.A0(\comb_reg_address[0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U128 (
	.Y(FE_OFN9_REG_ADDRESS_1_),
	.B1(n84),
	.B0(n29),
	.A1(n83),
	.A0(n99), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Reg_file_DATA_WIDTH8_ADDRESS_BITS3_test_1 (
	CLK, 
	RST, 
	R_REG_EN, 
	W_REG_EN, 
	REG_ADDRESS, 
	W_REG_DATA, 
	R_DATA_VALID, 
	R_REG_DATA, 
	REG0, 
	REG1, 
	REG2, 
	REG3, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN4_scanclkref, 
	FE_OFN5_scanclkref, 
	FE_OFN12_SE, 
	FE_OFN13_SE, 
	FE_OFN14_SE, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input R_REG_EN;
   input W_REG_EN;
   input [3:0] REG_ADDRESS;
   input [7:0] W_REG_DATA;
   output R_DATA_VALID;
   output [7:0] R_REG_DATA;
   output [7:0] REG0;
   output [7:0] REG1;
   output [7:0] REG2;
   output [7:0] REG3;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN4_scanclkref;
   input FE_OFN5_scanclkref;
   input FE_OFN12_SE;
   input FE_OFN13_SE;
   input FE_OFN14_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N10;
   wire N11;
   wire N12;
   wire N13;
   wire \Reg_file[15][7] ;
   wire \Reg_file[15][6] ;
   wire \Reg_file[15][5] ;
   wire \Reg_file[15][4] ;
   wire \Reg_file[15][3] ;
   wire \Reg_file[15][2] ;
   wire \Reg_file[15][1] ;
   wire \Reg_file[15][0] ;
   wire \Reg_file[14][7] ;
   wire \Reg_file[14][6] ;
   wire \Reg_file[14][5] ;
   wire \Reg_file[14][4] ;
   wire \Reg_file[14][3] ;
   wire \Reg_file[14][2] ;
   wire \Reg_file[14][1] ;
   wire \Reg_file[14][0] ;
   wire \Reg_file[13][7] ;
   wire \Reg_file[13][6] ;
   wire \Reg_file[13][5] ;
   wire \Reg_file[13][4] ;
   wire \Reg_file[13][3] ;
   wire \Reg_file[13][2] ;
   wire \Reg_file[13][1] ;
   wire \Reg_file[13][0] ;
   wire \Reg_file[12][7] ;
   wire \Reg_file[12][6] ;
   wire \Reg_file[12][5] ;
   wire \Reg_file[12][4] ;
   wire \Reg_file[12][3] ;
   wire \Reg_file[12][2] ;
   wire \Reg_file[12][1] ;
   wire \Reg_file[12][0] ;
   wire \Reg_file[11][7] ;
   wire \Reg_file[11][6] ;
   wire \Reg_file[11][5] ;
   wire \Reg_file[11][4] ;
   wire \Reg_file[11][3] ;
   wire \Reg_file[11][2] ;
   wire \Reg_file[11][1] ;
   wire \Reg_file[11][0] ;
   wire \Reg_file[10][7] ;
   wire \Reg_file[10][6] ;
   wire \Reg_file[10][5] ;
   wire \Reg_file[10][4] ;
   wire \Reg_file[10][3] ;
   wire \Reg_file[10][2] ;
   wire \Reg_file[10][1] ;
   wire \Reg_file[10][0] ;
   wire \Reg_file[9][7] ;
   wire \Reg_file[9][6] ;
   wire \Reg_file[9][5] ;
   wire \Reg_file[9][4] ;
   wire \Reg_file[9][3] ;
   wire \Reg_file[9][2] ;
   wire \Reg_file[9][1] ;
   wire \Reg_file[9][0] ;
   wire \Reg_file[8][7] ;
   wire \Reg_file[8][6] ;
   wire \Reg_file[8][5] ;
   wire \Reg_file[8][4] ;
   wire \Reg_file[8][3] ;
   wire \Reg_file[8][2] ;
   wire \Reg_file[8][1] ;
   wire \Reg_file[8][0] ;
   wire \Reg_file[7][7] ;
   wire \Reg_file[7][6] ;
   wire \Reg_file[7][5] ;
   wire \Reg_file[7][4] ;
   wire \Reg_file[7][3] ;
   wire \Reg_file[7][2] ;
   wire \Reg_file[7][1] ;
   wire \Reg_file[7][0] ;
   wire \Reg_file[6][7] ;
   wire \Reg_file[6][6] ;
   wire \Reg_file[6][5] ;
   wire \Reg_file[6][4] ;
   wire \Reg_file[6][3] ;
   wire \Reg_file[6][2] ;
   wire \Reg_file[6][1] ;
   wire \Reg_file[6][0] ;
   wire \Reg_file[5][7] ;
   wire \Reg_file[5][6] ;
   wire \Reg_file[5][5] ;
   wire \Reg_file[5][4] ;
   wire \Reg_file[5][3] ;
   wire \Reg_file[5][2] ;
   wire \Reg_file[5][1] ;
   wire \Reg_file[5][0] ;
   wire \Reg_file[4][7] ;
   wire \Reg_file[4][6] ;
   wire \Reg_file[4][5] ;
   wire \Reg_file[4][4] ;
   wire \Reg_file[4][3] ;
   wire \Reg_file[4][2] ;
   wire \Reg_file[4][1] ;
   wire \Reg_file[4][0] ;
   wire N35;
   wire N36;
   wire N37;
   wire N38;
   wire N39;
   wire N40;
   wire N41;
   wire N42;
   wire N59;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n336;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;

   assign N10 = REG_ADDRESS[0] ;
   assign N11 = REG_ADDRESS[1] ;
   assign N12 = REG_ADDRESS[2] ;
   assign N13 = REG_ADDRESS[3] ;
   assign test_so = \Reg_file[15][7]  ;

   // Module instantiations
   SDFFQX2M \R_REG_DATA_reg[7]  (
	.SI(R_REG_DATA[6]),
	.SE(test_se),
	.Q(R_REG_DATA[7]),
	.D(n185),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \R_REG_DATA_reg[6]  (
	.SI(R_REG_DATA[5]),
	.SE(test_se),
	.Q(R_REG_DATA[6]),
	.D(n184),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \R_REG_DATA_reg[5]  (
	.SI(R_REG_DATA[4]),
	.SE(test_se),
	.Q(R_REG_DATA[5]),
	.D(n183),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \R_REG_DATA_reg[4]  (
	.SI(R_REG_DATA[3]),
	.SE(test_se),
	.Q(R_REG_DATA[4]),
	.D(n182),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \R_REG_DATA_reg[3]  (
	.SI(R_REG_DATA[2]),
	.SE(test_se),
	.Q(R_REG_DATA[3]),
	.D(n181),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \R_REG_DATA_reg[2]  (
	.SI(R_REG_DATA[1]),
	.SE(test_se),
	.Q(R_REG_DATA[2]),
	.D(n180),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \R_REG_DATA_reg[1]  (
	.SI(R_REG_DATA[0]),
	.SE(test_se),
	.Q(R_REG_DATA[1]),
	.D(n179),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \R_REG_DATA_reg[0]  (
	.SI(R_DATA_VALID),
	.SE(test_se),
	.Q(R_REG_DATA[0]),
	.D(n178),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[13][7]  (
	.SI(\Reg_file[13][6] ),
	.SE(FE_OFN12_SE),
	.RN(n350),
	.Q(\Reg_file[13][7] ),
	.D(n297),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[13][6]  (
	.SI(\Reg_file[13][5] ),
	.SE(FE_OFN12_SE),
	.RN(n350),
	.Q(\Reg_file[13][6] ),
	.D(n296),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[13][5]  (
	.SI(\Reg_file[13][4] ),
	.SE(FE_OFN12_SE),
	.RN(n350),
	.Q(\Reg_file[13][5] ),
	.D(n295),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[13][4]  (
	.SI(\Reg_file[13][3] ),
	.SE(FE_OFN12_SE),
	.RN(n349),
	.Q(\Reg_file[13][4] ),
	.D(n294),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[13][3]  (
	.SI(\Reg_file[13][2] ),
	.SE(FE_OFN13_SE),
	.RN(n344),
	.Q(\Reg_file[13][3] ),
	.D(n293),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[13][2]  (
	.SI(\Reg_file[13][1] ),
	.SE(FE_OFN12_SE),
	.RN(n350),
	.Q(\Reg_file[13][2] ),
	.D(n292),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[13][1]  (
	.SI(\Reg_file[13][0] ),
	.SE(FE_OFN12_SE),
	.RN(n348),
	.Q(\Reg_file[13][1] ),
	.D(n291),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[13][0]  (
	.SI(\Reg_file[12][7] ),
	.SE(FE_OFN12_SE),
	.RN(n347),
	.Q(\Reg_file[13][0] ),
	.D(n290),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[9][7]  (
	.SI(\Reg_file[9][6] ),
	.SE(FE_OFN14_SE),
	.RN(n348),
	.Q(\Reg_file[9][7] ),
	.D(n265),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[9][6]  (
	.SI(\Reg_file[9][5] ),
	.SE(FE_OFN12_SE),
	.RN(n348),
	.Q(\Reg_file[9][6] ),
	.D(n264),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[9][5]  (
	.SI(\Reg_file[9][4] ),
	.SE(FE_OFN12_SE),
	.RN(n348),
	.Q(\Reg_file[9][5] ),
	.D(n263),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[9][4]  (
	.SI(\Reg_file[9][3] ),
	.SE(FE_OFN12_SE),
	.RN(n348),
	.Q(\Reg_file[9][4] ),
	.D(n262),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[9][3]  (
	.SI(\Reg_file[9][2] ),
	.SE(FE_OFN12_SE),
	.RN(n348),
	.Q(\Reg_file[9][3] ),
	.D(n261),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[9][2]  (
	.SI(\Reg_file[9][1] ),
	.SE(FE_OFN13_SE),
	.RN(n348),
	.Q(\Reg_file[9][2] ),
	.D(n260),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[9][1]  (
	.SI(\Reg_file[9][0] ),
	.SE(FE_OFN13_SE),
	.RN(n348),
	.Q(\Reg_file[9][1] ),
	.D(n259),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[9][0]  (
	.SI(\Reg_file[8][7] ),
	.SE(FE_OFN12_SE),
	.RN(n348),
	.Q(\Reg_file[9][0] ),
	.D(n258),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[5][7]  (
	.SI(\Reg_file[5][6] ),
	.SE(FE_OFN14_SE),
	.RN(n346),
	.Q(\Reg_file[5][7] ),
	.D(n233),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[5][6]  (
	.SI(\Reg_file[5][5] ),
	.SE(FE_OFN12_SE),
	.RN(n346),
	.Q(\Reg_file[5][6] ),
	.D(n232),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[5][5]  (
	.SI(\Reg_file[5][4] ),
	.SE(FE_OFN14_SE),
	.RN(n346),
	.Q(\Reg_file[5][5] ),
	.D(n231),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[5][4]  (
	.SI(\Reg_file[5][3] ),
	.SE(FE_OFN14_SE),
	.RN(n346),
	.Q(\Reg_file[5][4] ),
	.D(n230),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[5][3]  (
	.SI(\Reg_file[5][2] ),
	.SE(FE_OFN14_SE),
	.RN(n346),
	.Q(\Reg_file[5][3] ),
	.D(n229),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[5][2]  (
	.SI(\Reg_file[5][1] ),
	.SE(FE_OFN14_SE),
	.RN(n346),
	.Q(\Reg_file[5][2] ),
	.D(n228),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[5][1]  (
	.SI(\Reg_file[5][0] ),
	.SE(FE_OFN14_SE),
	.RN(n346),
	.Q(\Reg_file[5][1] ),
	.D(n227),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[5][0]  (
	.SI(\Reg_file[4][7] ),
	.SE(FE_OFN14_SE),
	.RN(n346),
	.Q(\Reg_file[5][0] ),
	.D(n226),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[15][7]  (
	.SI(\Reg_file[15][6] ),
	.SE(test_se),
	.RN(n344),
	.Q(\Reg_file[15][7] ),
	.D(n313),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[15][6]  (
	.SI(\Reg_file[15][5] ),
	.SE(FE_OFN12_SE),
	.RN(n345),
	.Q(\Reg_file[15][6] ),
	.D(n312),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[15][5]  (
	.SI(\Reg_file[15][4] ),
	.SE(FE_OFN12_SE),
	.RN(n348),
	.Q(\Reg_file[15][5] ),
	.D(n311),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[15][4]  (
	.SI(\Reg_file[15][3] ),
	.SE(FE_OFN12_SE),
	.RN(n347),
	.Q(\Reg_file[15][4] ),
	.D(n310),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[15][3]  (
	.SI(\Reg_file[15][2] ),
	.SE(FE_OFN13_SE),
	.RN(n346),
	.Q(\Reg_file[15][3] ),
	.D(n309),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[15][2]  (
	.SI(\Reg_file[15][1] ),
	.SE(FE_OFN13_SE),
	.RN(n350),
	.Q(\Reg_file[15][2] ),
	.D(n308),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[15][1]  (
	.SI(\Reg_file[15][0] ),
	.SE(FE_OFN13_SE),
	.RN(n350),
	.Q(\Reg_file[15][1] ),
	.D(n307),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[15][0]  (
	.SI(\Reg_file[14][7] ),
	.SE(FE_OFN12_SE),
	.RN(n350),
	.Q(\Reg_file[15][0] ),
	.D(n306),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[11][7]  (
	.SI(\Reg_file[11][6] ),
	.SE(FE_OFN12_SE),
	.RN(n346),
	.Q(\Reg_file[11][7] ),
	.D(n281),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[11][6]  (
	.SI(\Reg_file[11][5] ),
	.SE(FE_OFN14_SE),
	.RN(n349),
	.Q(\Reg_file[11][6] ),
	.D(n280),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[11][5]  (
	.SI(\Reg_file[11][4] ),
	.SE(FE_OFN12_SE),
	.RN(n349),
	.Q(\Reg_file[11][5] ),
	.D(n279),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[11][4]  (
	.SI(\Reg_file[11][3] ),
	.SE(FE_OFN12_SE),
	.RN(n349),
	.Q(\Reg_file[11][4] ),
	.D(n278),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[11][3]  (
	.SI(\Reg_file[11][2] ),
	.SE(FE_OFN12_SE),
	.RN(n349),
	.Q(\Reg_file[11][3] ),
	.D(n277),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[11][2]  (
	.SI(\Reg_file[11][1] ),
	.SE(FE_OFN12_SE),
	.RN(n349),
	.Q(\Reg_file[11][2] ),
	.D(n276),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[11][1]  (
	.SI(\Reg_file[11][0] ),
	.SE(FE_OFN12_SE),
	.RN(n349),
	.Q(\Reg_file[11][1] ),
	.D(n275),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[11][0]  (
	.SI(\Reg_file[10][7] ),
	.SE(FE_OFN12_SE),
	.RN(n349),
	.Q(\Reg_file[11][0] ),
	.D(n274),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[7][7]  (
	.SI(\Reg_file[7][6] ),
	.SE(FE_OFN14_SE),
	.RN(n347),
	.Q(\Reg_file[7][7] ),
	.D(n249),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[7][6]  (
	.SI(\Reg_file[7][5] ),
	.SE(FE_OFN14_SE),
	.RN(n347),
	.Q(\Reg_file[7][6] ),
	.D(n248),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[7][5]  (
	.SI(\Reg_file[7][4] ),
	.SE(FE_OFN14_SE),
	.RN(n347),
	.Q(\Reg_file[7][5] ),
	.D(n247),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[7][4]  (
	.SI(\Reg_file[7][3] ),
	.SE(FE_OFN14_SE),
	.RN(n347),
	.Q(\Reg_file[7][4] ),
	.D(n246),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[7][3]  (
	.SI(\Reg_file[7][2] ),
	.SE(FE_OFN14_SE),
	.RN(n347),
	.Q(\Reg_file[7][3] ),
	.D(n245),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[7][2]  (
	.SI(\Reg_file[7][1] ),
	.SE(FE_OFN14_SE),
	.RN(n347),
	.Q(\Reg_file[7][2] ),
	.D(n244),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[7][1]  (
	.SI(\Reg_file[7][0] ),
	.SE(FE_OFN14_SE),
	.RN(n347),
	.Q(\Reg_file[7][1] ),
	.D(n243),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[7][0]  (
	.SI(\Reg_file[6][7] ),
	.SE(FE_OFN14_SE),
	.RN(n347),
	.Q(\Reg_file[7][0] ),
	.D(n242),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[14][7]  (
	.SI(\Reg_file[14][6] ),
	.SE(FE_OFN12_SE),
	.RN(n350),
	.Q(\Reg_file[14][7] ),
	.D(n305),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[14][6]  (
	.SI(\Reg_file[14][5] ),
	.SE(FE_OFN12_SE),
	.RN(n350),
	.Q(\Reg_file[14][6] ),
	.D(n304),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[14][5]  (
	.SI(\Reg_file[14][4] ),
	.SE(FE_OFN12_SE),
	.RN(n350),
	.Q(\Reg_file[14][5] ),
	.D(n303),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[14][4]  (
	.SI(\Reg_file[14][3] ),
	.SE(FE_OFN12_SE),
	.RN(n350),
	.Q(\Reg_file[14][4] ),
	.D(n302),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[14][3]  (
	.SI(\Reg_file[14][2] ),
	.SE(FE_OFN12_SE),
	.RN(n350),
	.Q(\Reg_file[14][3] ),
	.D(n301),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[14][2]  (
	.SI(\Reg_file[14][1] ),
	.SE(FE_OFN12_SE),
	.RN(n350),
	.Q(\Reg_file[14][2] ),
	.D(n300),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[14][1]  (
	.SI(\Reg_file[14][0] ),
	.SE(FE_OFN12_SE),
	.RN(n350),
	.Q(\Reg_file[14][1] ),
	.D(n299),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[14][0]  (
	.SI(\Reg_file[13][7] ),
	.SE(FE_OFN12_SE),
	.RN(n350),
	.Q(\Reg_file[14][0] ),
	.D(n298),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[10][7]  (
	.SI(\Reg_file[10][6] ),
	.SE(FE_OFN14_SE),
	.RN(n349),
	.Q(\Reg_file[10][7] ),
	.D(n273),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[10][6]  (
	.SI(\Reg_file[10][5] ),
	.SE(FE_OFN14_SE),
	.RN(n349),
	.Q(\Reg_file[10][6] ),
	.D(n272),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[10][5]  (
	.SI(\Reg_file[10][4] ),
	.SE(FE_OFN12_SE),
	.RN(n349),
	.Q(\Reg_file[10][5] ),
	.D(n271),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[10][4]  (
	.SI(\Reg_file[10][3] ),
	.SE(FE_OFN12_SE),
	.RN(n349),
	.Q(\Reg_file[10][4] ),
	.D(n270),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[10][3]  (
	.SI(\Reg_file[10][2] ),
	.SE(FE_OFN12_SE),
	.RN(n349),
	.Q(\Reg_file[10][3] ),
	.D(n269),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[10][2]  (
	.SI(\Reg_file[10][1] ),
	.SE(FE_OFN13_SE),
	.RN(n349),
	.Q(\Reg_file[10][2] ),
	.D(n268),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[10][1]  (
	.SI(\Reg_file[10][0] ),
	.SE(FE_OFN13_SE),
	.RN(n349),
	.Q(\Reg_file[10][1] ),
	.D(n267),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[10][0]  (
	.SI(\Reg_file[9][7] ),
	.SE(FE_OFN12_SE),
	.RN(n348),
	.Q(\Reg_file[10][0] ),
	.D(n266),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[6][7]  (
	.SI(\Reg_file[6][6] ),
	.SE(FE_OFN14_SE),
	.RN(n347),
	.Q(\Reg_file[6][7] ),
	.D(n241),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[6][6]  (
	.SI(\Reg_file[6][5] ),
	.SE(FE_OFN12_SE),
	.RN(n347),
	.Q(\Reg_file[6][6] ),
	.D(n240),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[6][5]  (
	.SI(\Reg_file[6][4] ),
	.SE(FE_OFN12_SE),
	.RN(n346),
	.Q(\Reg_file[6][5] ),
	.D(n239),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[6][4]  (
	.SI(\Reg_file[6][3] ),
	.SE(FE_OFN14_SE),
	.RN(n346),
	.Q(\Reg_file[6][4] ),
	.D(n238),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[6][3]  (
	.SI(\Reg_file[6][2] ),
	.SE(FE_OFN14_SE),
	.RN(n346),
	.Q(\Reg_file[6][3] ),
	.D(n237),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[6][2]  (
	.SI(\Reg_file[6][1] ),
	.SE(FE_OFN14_SE),
	.RN(n346),
	.Q(\Reg_file[6][2] ),
	.D(n236),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[6][1]  (
	.SI(\Reg_file[6][0] ),
	.SE(FE_OFN14_SE),
	.RN(n346),
	.Q(\Reg_file[6][1] ),
	.D(n235),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[6][0]  (
	.SI(\Reg_file[5][7] ),
	.SE(FE_OFN14_SE),
	.RN(n346),
	.Q(\Reg_file[6][0] ),
	.D(n234),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[12][7]  (
	.SI(\Reg_file[12][6] ),
	.SE(FE_OFN12_SE),
	.RN(n345),
	.Q(\Reg_file[12][7] ),
	.D(n289),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[12][6]  (
	.SI(\Reg_file[12][5] ),
	.SE(FE_OFN12_SE),
	.RN(n345),
	.Q(\Reg_file[12][6] ),
	.D(n288),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[12][5]  (
	.SI(\Reg_file[12][4] ),
	.SE(FE_OFN12_SE),
	.RN(n349),
	.Q(\Reg_file[12][5] ),
	.D(n287),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[12][4]  (
	.SI(\Reg_file[12][3] ),
	.SE(FE_OFN12_SE),
	.RN(n344),
	.Q(\Reg_file[12][4] ),
	.D(n286),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[12][3]  (
	.SI(\Reg_file[12][2] ),
	.SE(FE_OFN13_SE),
	.RN(n350),
	.Q(\Reg_file[12][3] ),
	.D(n285),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[12][2]  (
	.SI(\Reg_file[12][1] ),
	.SE(FE_OFN13_SE),
	.RN(n348),
	.Q(\Reg_file[12][2] ),
	.D(n284),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[12][1]  (
	.SI(\Reg_file[12][0] ),
	.SE(FE_OFN13_SE),
	.RN(n347),
	.Q(\Reg_file[12][1] ),
	.D(n283),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[12][0]  (
	.SI(\Reg_file[11][7] ),
	.SE(FE_OFN12_SE),
	.RN(n346),
	.Q(\Reg_file[12][0] ),
	.D(n282),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[8][7]  (
	.SI(\Reg_file[8][6] ),
	.SE(FE_OFN12_SE),
	.RN(n348),
	.Q(\Reg_file[8][7] ),
	.D(n257),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[8][6]  (
	.SI(\Reg_file[8][5] ),
	.SE(FE_OFN12_SE),
	.RN(n348),
	.Q(\Reg_file[8][6] ),
	.D(n256),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[8][5]  (
	.SI(\Reg_file[8][4] ),
	.SE(FE_OFN12_SE),
	.RN(n348),
	.Q(\Reg_file[8][5] ),
	.D(n255),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[8][4]  (
	.SI(\Reg_file[8][3] ),
	.SE(FE_OFN12_SE),
	.RN(n348),
	.Q(\Reg_file[8][4] ),
	.D(n254),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[8][3]  (
	.SI(\Reg_file[8][2] ),
	.SE(FE_OFN12_SE),
	.RN(n348),
	.Q(\Reg_file[8][3] ),
	.D(n253),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[8][2]  (
	.SI(\Reg_file[8][1] ),
	.SE(FE_OFN12_SE),
	.RN(n347),
	.Q(\Reg_file[8][2] ),
	.D(n252),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[8][1]  (
	.SI(\Reg_file[8][0] ),
	.SE(FE_OFN12_SE),
	.RN(n347),
	.Q(\Reg_file[8][1] ),
	.D(n251),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[8][0]  (
	.SI(\Reg_file[7][7] ),
	.SE(FE_OFN14_SE),
	.RN(n347),
	.Q(\Reg_file[8][0] ),
	.D(n250),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[4][7]  (
	.SI(\Reg_file[4][6] ),
	.SE(FE_OFN14_SE),
	.RN(n345),
	.Q(\Reg_file[4][7] ),
	.D(n225),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[4][6]  (
	.SI(\Reg_file[4][5] ),
	.SE(FE_OFN14_SE),
	.RN(n345),
	.Q(\Reg_file[4][6] ),
	.D(n224),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[4][5]  (
	.SI(\Reg_file[4][4] ),
	.SE(FE_OFN14_SE),
	.RN(n345),
	.Q(\Reg_file[4][5] ),
	.D(n223),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[4][4]  (
	.SI(\Reg_file[4][3] ),
	.SE(FE_OFN14_SE),
	.RN(n345),
	.Q(\Reg_file[4][4] ),
	.D(n222),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[4][3]  (
	.SI(\Reg_file[4][2] ),
	.SE(FE_OFN14_SE),
	.RN(n345),
	.Q(\Reg_file[4][3] ),
	.D(n221),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[4][2]  (
	.SI(\Reg_file[4][1] ),
	.SE(FE_OFN14_SE),
	.RN(n345),
	.Q(\Reg_file[4][2] ),
	.D(n220),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[4][1]  (
	.SI(\Reg_file[4][0] ),
	.SE(test_se),
	.RN(n345),
	.Q(\Reg_file[4][1] ),
	.D(n219),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[4][0]  (
	.SI(REG3[7]),
	.SE(test_se),
	.RN(n345),
	.Q(\Reg_file[4][0] ),
	.D(n218),
	.CK(FE_OFN4_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[3][0]  (
	.SI(REG2[7]),
	.SE(test_se),
	.RN(n344),
	.Q(REG3[0]),
	.D(n210),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[2][1]  (
	.SI(REG2[0]),
	.SE(test_se),
	.RN(n344),
	.Q(REG2[1]),
	.D(n203),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[1][6]  (
	.SI(REG1[5]),
	.SE(test_se),
	.RN(n344),
	.Q(REG1[6]),
	.D(n200),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[0][7]  (
	.SI(REG0[6]),
	.SE(test_se),
	.RN(n349),
	.Q(REG0[7]),
	.D(n193),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[0][6]  (
	.SI(REG0[5]),
	.SE(test_se),
	.RN(n350),
	.Q(REG0[6]),
	.D(n192),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[0][5]  (
	.SI(REG0[4]),
	.SE(test_se),
	.RN(n348),
	.Q(REG0[5]),
	.D(n191),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[0][4]  (
	.SI(REG0[3]),
	.SE(test_se),
	.RN(n347),
	.Q(REG0[4]),
	.D(n190),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[0][3]  (
	.SI(REG0[2]),
	.SE(test_se),
	.RN(n346),
	.Q(REG0[3]),
	.D(n189),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[0][2]  (
	.SI(REG0[1]),
	.SE(test_se),
	.RN(n345),
	.Q(REG0[2]),
	.D(n188),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[0][1]  (
	.SI(REG0[0]),
	.SE(test_se),
	.RN(n344),
	.Q(REG0[1]),
	.D(n187),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[0][0]  (
	.SI(R_REG_DATA[7]),
	.SE(test_se),
	.RN(n349),
	.Q(REG0[0]),
	.D(n186),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M R_DATA_VALID_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(n347),
	.Q(R_DATA_VALID),
	.D(N59),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \Reg_file_reg[3][5]  (
	.SN(n347),
	.SI(REG3[4]),
	.SE(test_se),
	.Q(REG3[5]),
	.D(n215),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[3][1]  (
	.SI(REG3[0]),
	.SE(test_se),
	.RN(n345),
	.Q(REG3[1]),
	.D(n211),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[3][4]  (
	.SI(REG3[3]),
	.SE(test_se),
	.RN(n345),
	.Q(REG3[4]),
	.D(n214),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[3][6]  (
	.SI(REG3[5]),
	.SE(test_se),
	.RN(n345),
	.Q(REG3[6]),
	.D(n216),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[3][3]  (
	.SI(REG3[2]),
	.SE(test_se),
	.RN(n345),
	.Q(REG3[3]),
	.D(n213),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[3][2]  (
	.SI(REG3[1]),
	.SE(test_se),
	.RN(n345),
	.Q(REG3[2]),
	.D(n212),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[3][7]  (
	.SI(REG3[6]),
	.SE(test_se),
	.RN(n345),
	.Q(REG3[7]),
	.D(n217),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \Reg_file_reg[2][0]  (
	.SN(n346),
	.SI(REG1[7]),
	.SE(test_se),
	.Q(REG2[0]),
	.D(n202),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[2][4]  (
	.SI(REG2[3]),
	.SE(test_se),
	.RN(n344),
	.Q(REG2[4]),
	.D(n206),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[2][2]  (
	.SI(REG2[1]),
	.SE(test_se),
	.RN(n344),
	.Q(REG2[2]),
	.D(n204),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[1][1]  (
	.SI(REG1[0]),
	.SE(test_se),
	.RN(n350),
	.Q(REG1[1]),
	.D(n195),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[1][5]  (
	.SI(REG1[4]),
	.SE(test_se),
	.RN(n344),
	.Q(REG1[5]),
	.D(n199),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[1][4]  (
	.SI(REG1[3]),
	.SE(test_se),
	.RN(n344),
	.Q(REG1[4]),
	.D(n198),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[1][7]  (
	.SI(REG1[6]),
	.SE(test_se),
	.RN(n344),
	.Q(REG1[7]),
	.D(n201),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \Reg_file_reg[2][7]  (
	.SN(n345),
	.SI(REG2[6]),
	.SE(test_se),
	.Q(REG2[7]),
	.D(n209),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[2][3]  (
	.SI(REG2[2]),
	.SE(test_se),
	.RN(n344),
	.Q(REG2[3]),
	.D(n205),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[1][3]  (
	.SI(REG1[2]),
	.SE(test_se),
	.RN(n344),
	.Q(REG1[3]),
	.D(n197),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[1][2]  (
	.SI(REG1[1]),
	.SE(test_se),
	.RN(n344),
	.Q(REG1[2]),
	.D(n196),
	.CK(FE_OFN5_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[2][5]  (
	.SI(REG2[4]),
	.SE(test_se),
	.RN(n344),
	.Q(REG2[5]),
	.D(n207),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[2][6]  (
	.SI(REG2[5]),
	.SE(test_se),
	.RN(n344),
	.Q(REG2[6]),
	.D(n208),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_file_reg[1][0]  (
	.SI(REG0[7]),
	.SE(test_se),
	.RN(n344),
	.Q(REG1[0]),
	.D(n194),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U140 (
	.Y(n170),
	.B(n341),
	.AN(n176), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U141 (
	.Y(n161),
	.B(N11),
	.AN(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U142 (
	.Y(n164),
	.B(n342),
	.AN(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U143 (
	.Y(n158),
	.B(N12),
	.A(n342), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U144 (
	.Y(n153),
	.B(N12),
	.A(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U145 (
	.Y(n156),
	.B(n341),
	.AN(n165), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U146 (
	.Y(n339),
	.A(n341), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U147 (
	.Y(n338),
	.A(n341), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U148 (
	.Y(n336),
	.A(n342), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U149 (
	.Y(n350),
	.A(n343), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U150 (
	.Y(n344),
	.A(n343), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U151 (
	.Y(n345),
	.A(n343), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX4M U152 (
	.Y(n346),
	.A(n343), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX4M U153 (
	.Y(n347),
	.A(n343), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U154 (
	.Y(n348),
	.A(n343), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U155 (
	.Y(n349),
	.A(n343), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U156 (
	.Y(n150),
	.B(n149),
	.AN(N59), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U157 (
	.Y(n149),
	.B(n343),
	.A(n151), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U158 (
	.Y(n340),
	.A(n341), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U166 (
	.Y(n154),
	.B(N10),
	.AN(n165), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U167 (
	.Y(n168),
	.B(N10),
	.AN(n176), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U168 (
	.Y(n155),
	.B(n153),
	.A(n156), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U169 (
	.Y(n167),
	.B(n153),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U170 (
	.Y(n169),
	.B(n153),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U171 (
	.Y(n171),
	.B(n158),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U172 (
	.Y(n172),
	.B(n158),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U173 (
	.Y(n157),
	.B(n154),
	.A(n158), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U174 (
	.Y(n159),
	.B(n156),
	.A(n158), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U175 (
	.Y(n160),
	.B(n154),
	.A(n161), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U176 (
	.Y(n162),
	.B(n156),
	.A(n161), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U177 (
	.Y(n163),
	.B(n154),
	.A(n164), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U178 (
	.Y(n166),
	.B(n156),
	.A(n164), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U179 (
	.Y(n173),
	.B(n161),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U180 (
	.Y(n174),
	.B(n161),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U181 (
	.Y(n175),
	.B(n164),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U182 (
	.Y(n177),
	.B(n164),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U183 (
	.Y(n152),
	.B(n154),
	.A(n153), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U184 (
	.Y(n151),
	.B(R_REG_EN),
	.AN(W_REG_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U185 (
	.Y(N59),
	.B(W_REG_EN),
	.AN(R_REG_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U192 (
	.Y(n366),
	.A(W_REG_DATA[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U193 (
	.Y(n368),
	.A(W_REG_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U194 (
	.Y(n369),
	.A(W_REG_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U195 (
	.Y(n370),
	.A(W_REG_DATA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U196 (
	.Y(n371),
	.A(W_REG_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U197 (
	.Y(n372),
	.A(W_REG_DATA[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U198 (
	.Y(n373),
	.A(W_REG_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U199 (
	.Y(n367),
	.A(W_REG_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U200 (
	.Y(n165),
	.B(N13),
	.AN(n151), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U201 (
	.Y(n176),
	.B(n151),
	.A(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U206 (
	.Y(n343),
	.A(RST), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U207 (
	.Y(n186),
	.B1(n366),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U208 (
	.Y(n187),
	.B1(n367),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U209 (
	.Y(n188),
	.B1(n368),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U210 (
	.Y(n189),
	.B1(n369),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U211 (
	.Y(n190),
	.B1(n370),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U212 (
	.Y(n191),
	.B1(n371),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U213 (
	.Y(n192),
	.B1(n372),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U214 (
	.Y(n193),
	.B1(n373),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U215 (
	.Y(n194),
	.B1(n155),
	.B0(n366),
	.A1N(n155),
	.A0N(REG1[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U216 (
	.Y(n195),
	.B1(n155),
	.B0(n367),
	.A1N(n155),
	.A0N(REG1[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U217 (
	.Y(n196),
	.B1(n155),
	.B0(n368),
	.A1N(n155),
	.A0N(REG1[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U218 (
	.Y(n197),
	.B1(n155),
	.B0(n369),
	.A1N(n155),
	.A0N(REG1[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U219 (
	.Y(n198),
	.B1(n155),
	.B0(n370),
	.A1N(n155),
	.A0N(REG1[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U220 (
	.Y(n199),
	.B1(n155),
	.B0(n371),
	.A1N(n155),
	.A0N(REG1[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U221 (
	.Y(n200),
	.B1(n155),
	.B0(n372),
	.A1N(n155),
	.A0N(REG1[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U222 (
	.Y(n201),
	.B1(n155),
	.B0(n373),
	.A1N(n155),
	.A0N(REG1[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U223 (
	.Y(n218),
	.B1(n160),
	.B0(n366),
	.A1N(n160),
	.A0N(\Reg_file[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U224 (
	.Y(n219),
	.B1(n160),
	.B0(n367),
	.A1N(n160),
	.A0N(\Reg_file[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U225 (
	.Y(n220),
	.B1(n160),
	.B0(n368),
	.A1N(n160),
	.A0N(\Reg_file[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U226 (
	.Y(n221),
	.B1(n160),
	.B0(n369),
	.A1N(n160),
	.A0N(\Reg_file[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U227 (
	.Y(n222),
	.B1(n160),
	.B0(n370),
	.A1N(n160),
	.A0N(\Reg_file[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U228 (
	.Y(n223),
	.B1(n160),
	.B0(n371),
	.A1N(n160),
	.A0N(\Reg_file[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U229 (
	.Y(n224),
	.B1(n160),
	.B0(n372),
	.A1N(n160),
	.A0N(\Reg_file[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U230 (
	.Y(n225),
	.B1(n160),
	.B0(n373),
	.A1N(n160),
	.A0N(\Reg_file[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U231 (
	.Y(n226),
	.B1(n162),
	.B0(n366),
	.A1N(n162),
	.A0N(\Reg_file[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U232 (
	.Y(n227),
	.B1(n162),
	.B0(n367),
	.A1N(n162),
	.A0N(\Reg_file[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U233 (
	.Y(n228),
	.B1(n162),
	.B0(n368),
	.A1N(n162),
	.A0N(\Reg_file[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U234 (
	.Y(n229),
	.B1(n162),
	.B0(n369),
	.A1N(n162),
	.A0N(\Reg_file[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U235 (
	.Y(n230),
	.B1(n162),
	.B0(n370),
	.A1N(n162),
	.A0N(\Reg_file[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U236 (
	.Y(n231),
	.B1(n162),
	.B0(n371),
	.A1N(n162),
	.A0N(\Reg_file[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U237 (
	.Y(n232),
	.B1(n162),
	.B0(n372),
	.A1N(n162),
	.A0N(\Reg_file[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U238 (
	.Y(n233),
	.B1(n162),
	.B0(n373),
	.A1N(n162),
	.A0N(\Reg_file[5][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U239 (
	.Y(n234),
	.B1(n163),
	.B0(n366),
	.A1N(n163),
	.A0N(\Reg_file[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U240 (
	.Y(n235),
	.B1(n163),
	.B0(n367),
	.A1N(n163),
	.A0N(\Reg_file[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U241 (
	.Y(n236),
	.B1(n163),
	.B0(n368),
	.A1N(n163),
	.A0N(\Reg_file[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U242 (
	.Y(n237),
	.B1(n163),
	.B0(n369),
	.A1N(n163),
	.A0N(\Reg_file[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U243 (
	.Y(n238),
	.B1(n163),
	.B0(n370),
	.A1N(n163),
	.A0N(\Reg_file[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U244 (
	.Y(n239),
	.B1(n163),
	.B0(n371),
	.A1N(n163),
	.A0N(\Reg_file[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U245 (
	.Y(n240),
	.B1(n163),
	.B0(n372),
	.A1N(n163),
	.A0N(\Reg_file[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U246 (
	.Y(n241),
	.B1(n163),
	.B0(n373),
	.A1N(n163),
	.A0N(\Reg_file[6][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U247 (
	.Y(n242),
	.B1(n166),
	.B0(n366),
	.A1N(n166),
	.A0N(\Reg_file[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U248 (
	.Y(n243),
	.B1(n166),
	.B0(n367),
	.A1N(n166),
	.A0N(\Reg_file[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U249 (
	.Y(n244),
	.B1(n166),
	.B0(n368),
	.A1N(n166),
	.A0N(\Reg_file[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U250 (
	.Y(n245),
	.B1(n166),
	.B0(n369),
	.A1N(n166),
	.A0N(\Reg_file[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U251 (
	.Y(n246),
	.B1(n166),
	.B0(n370),
	.A1N(n166),
	.A0N(\Reg_file[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U252 (
	.Y(n247),
	.B1(n166),
	.B0(n371),
	.A1N(n166),
	.A0N(\Reg_file[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U253 (
	.Y(n248),
	.B1(n166),
	.B0(n372),
	.A1N(n166),
	.A0N(\Reg_file[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U254 (
	.Y(n249),
	.B1(n166),
	.B0(n373),
	.A1N(n166),
	.A0N(\Reg_file[7][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U255 (
	.Y(n250),
	.B1(n167),
	.B0(n366),
	.A1N(n167),
	.A0N(\Reg_file[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U256 (
	.Y(n251),
	.B1(n167),
	.B0(n367),
	.A1N(n167),
	.A0N(\Reg_file[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U257 (
	.Y(n252),
	.B1(n167),
	.B0(n368),
	.A1N(n167),
	.A0N(\Reg_file[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U258 (
	.Y(n253),
	.B1(n167),
	.B0(n369),
	.A1N(n167),
	.A0N(\Reg_file[8][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U259 (
	.Y(n254),
	.B1(n167),
	.B0(n370),
	.A1N(n167),
	.A0N(\Reg_file[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U260 (
	.Y(n255),
	.B1(n167),
	.B0(n371),
	.A1N(n167),
	.A0N(\Reg_file[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U261 (
	.Y(n256),
	.B1(n167),
	.B0(n372),
	.A1N(n167),
	.A0N(\Reg_file[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U262 (
	.Y(n257),
	.B1(n167),
	.B0(n373),
	.A1N(n167),
	.A0N(\Reg_file[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U263 (
	.Y(n258),
	.B1(n169),
	.B0(n366),
	.A1N(n169),
	.A0N(\Reg_file[9][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U264 (
	.Y(n259),
	.B1(n169),
	.B0(n367),
	.A1N(n169),
	.A0N(\Reg_file[9][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U265 (
	.Y(n260),
	.B1(n169),
	.B0(n368),
	.A1N(n169),
	.A0N(\Reg_file[9][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U266 (
	.Y(n261),
	.B1(n169),
	.B0(n369),
	.A1N(n169),
	.A0N(\Reg_file[9][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U267 (
	.Y(n262),
	.B1(n169),
	.B0(n370),
	.A1N(n169),
	.A0N(\Reg_file[9][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U268 (
	.Y(n263),
	.B1(n169),
	.B0(n371),
	.A1N(n169),
	.A0N(\Reg_file[9][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U269 (
	.Y(n264),
	.B1(n169),
	.B0(n372),
	.A1N(n169),
	.A0N(\Reg_file[9][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U270 (
	.Y(n265),
	.B1(n169),
	.B0(n373),
	.A1N(n169),
	.A0N(\Reg_file[9][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U271 (
	.Y(n266),
	.B1(n171),
	.B0(n366),
	.A1N(n171),
	.A0N(\Reg_file[10][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U272 (
	.Y(n267),
	.B1(n171),
	.B0(n367),
	.A1N(n171),
	.A0N(\Reg_file[10][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U273 (
	.Y(n268),
	.B1(n171),
	.B0(n368),
	.A1N(n171),
	.A0N(\Reg_file[10][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U274 (
	.Y(n269),
	.B1(n171),
	.B0(n369),
	.A1N(n171),
	.A0N(\Reg_file[10][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U275 (
	.Y(n270),
	.B1(n171),
	.B0(n370),
	.A1N(n171),
	.A0N(\Reg_file[10][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U276 (
	.Y(n271),
	.B1(n171),
	.B0(n371),
	.A1N(n171),
	.A0N(\Reg_file[10][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U277 (
	.Y(n272),
	.B1(n171),
	.B0(n372),
	.A1N(n171),
	.A0N(\Reg_file[10][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U278 (
	.Y(n273),
	.B1(n171),
	.B0(n373),
	.A1N(n171),
	.A0N(\Reg_file[10][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U279 (
	.Y(n274),
	.B1(n172),
	.B0(n366),
	.A1N(n172),
	.A0N(\Reg_file[11][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U280 (
	.Y(n275),
	.B1(n172),
	.B0(n367),
	.A1N(n172),
	.A0N(\Reg_file[11][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U281 (
	.Y(n276),
	.B1(n172),
	.B0(n368),
	.A1N(n172),
	.A0N(\Reg_file[11][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U282 (
	.Y(n277),
	.B1(n172),
	.B0(n369),
	.A1N(n172),
	.A0N(\Reg_file[11][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U283 (
	.Y(n278),
	.B1(n172),
	.B0(n370),
	.A1N(n172),
	.A0N(\Reg_file[11][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U284 (
	.Y(n279),
	.B1(n172),
	.B0(n371),
	.A1N(n172),
	.A0N(\Reg_file[11][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U285 (
	.Y(n280),
	.B1(n172),
	.B0(n372),
	.A1N(n172),
	.A0N(\Reg_file[11][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U286 (
	.Y(n281),
	.B1(n172),
	.B0(n373),
	.A1N(n172),
	.A0N(\Reg_file[11][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U287 (
	.Y(n282),
	.B1(n173),
	.B0(n366),
	.A1N(n173),
	.A0N(\Reg_file[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U288 (
	.Y(n283),
	.B1(n173),
	.B0(n367),
	.A1N(n173),
	.A0N(\Reg_file[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U289 (
	.Y(n284),
	.B1(n173),
	.B0(n368),
	.A1N(n173),
	.A0N(\Reg_file[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U290 (
	.Y(n285),
	.B1(n173),
	.B0(n369),
	.A1N(n173),
	.A0N(\Reg_file[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U291 (
	.Y(n286),
	.B1(n173),
	.B0(n370),
	.A1N(n173),
	.A0N(\Reg_file[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U292 (
	.Y(n287),
	.B1(n173),
	.B0(n371),
	.A1N(n173),
	.A0N(\Reg_file[12][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U293 (
	.Y(n288),
	.B1(n173),
	.B0(n372),
	.A1N(n173),
	.A0N(\Reg_file[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U294 (
	.Y(n289),
	.B1(n173),
	.B0(n373),
	.A1N(n173),
	.A0N(\Reg_file[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U295 (
	.Y(n290),
	.B1(n174),
	.B0(n366),
	.A1N(n174),
	.A0N(\Reg_file[13][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U296 (
	.Y(n291),
	.B1(n174),
	.B0(n367),
	.A1N(n174),
	.A0N(\Reg_file[13][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U297 (
	.Y(n292),
	.B1(n174),
	.B0(n368),
	.A1N(n174),
	.A0N(\Reg_file[13][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U298 (
	.Y(n293),
	.B1(n174),
	.B0(n369),
	.A1N(n174),
	.A0N(\Reg_file[13][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U299 (
	.Y(n294),
	.B1(n174),
	.B0(n370),
	.A1N(n174),
	.A0N(\Reg_file[13][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U300 (
	.Y(n295),
	.B1(n174),
	.B0(n371),
	.A1N(n174),
	.A0N(\Reg_file[13][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U301 (
	.Y(n296),
	.B1(n174),
	.B0(n372),
	.A1N(n174),
	.A0N(\Reg_file[13][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U302 (
	.Y(n297),
	.B1(n174),
	.B0(n373),
	.A1N(n174),
	.A0N(\Reg_file[13][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U303 (
	.Y(n298),
	.B1(n175),
	.B0(n366),
	.A1N(n175),
	.A0N(\Reg_file[14][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U304 (
	.Y(n299),
	.B1(n175),
	.B0(n367),
	.A1N(n175),
	.A0N(\Reg_file[14][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U305 (
	.Y(n300),
	.B1(n175),
	.B0(n368),
	.A1N(n175),
	.A0N(\Reg_file[14][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U306 (
	.Y(n301),
	.B1(n175),
	.B0(n369),
	.A1N(n175),
	.A0N(\Reg_file[14][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U307 (
	.Y(n302),
	.B1(n175),
	.B0(n370),
	.A1N(n175),
	.A0N(\Reg_file[14][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U308 (
	.Y(n303),
	.B1(n175),
	.B0(n371),
	.A1N(n175),
	.A0N(\Reg_file[14][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U309 (
	.Y(n304),
	.B1(n175),
	.B0(n372),
	.A1N(n175),
	.A0N(\Reg_file[14][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U310 (
	.Y(n305),
	.B1(n175),
	.B0(n373),
	.A1N(n175),
	.A0N(\Reg_file[14][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U311 (
	.Y(n306),
	.B1(n177),
	.B0(n366),
	.A1N(n177),
	.A0N(\Reg_file[15][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U312 (
	.Y(n307),
	.B1(n177),
	.B0(n367),
	.A1N(n177),
	.A0N(\Reg_file[15][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U313 (
	.Y(n308),
	.B1(n177),
	.B0(n368),
	.A1N(n177),
	.A0N(\Reg_file[15][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U314 (
	.Y(n309),
	.B1(n177),
	.B0(n369),
	.A1N(n177),
	.A0N(\Reg_file[15][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U315 (
	.Y(n310),
	.B1(n177),
	.B0(n370),
	.A1N(n177),
	.A0N(\Reg_file[15][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U316 (
	.Y(n311),
	.B1(n177),
	.B0(n371),
	.A1N(n177),
	.A0N(\Reg_file[15][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U317 (
	.Y(n312),
	.B1(n177),
	.B0(n372),
	.A1N(n177),
	.A0N(\Reg_file[15][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U318 (
	.Y(n313),
	.B1(n177),
	.B0(n373),
	.A1N(n177),
	.A0N(\Reg_file[15][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U319 (
	.Y(n203),
	.B1(n157),
	.B0(n367),
	.A1N(n157),
	.A0N(REG2[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U320 (
	.Y(n204),
	.B1(n157),
	.B0(n368),
	.A1N(n157),
	.A0N(REG2[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U321 (
	.Y(n205),
	.B1(n157),
	.B0(n369),
	.A1N(n157),
	.A0N(REG2[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U322 (
	.Y(n206),
	.B1(n157),
	.B0(n370),
	.A1N(n157),
	.A0N(REG2[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U323 (
	.Y(n207),
	.B1(n157),
	.B0(n371),
	.A1N(n157),
	.A0N(REG2[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U324 (
	.Y(n208),
	.B1(n157),
	.B0(n372),
	.A1N(n157),
	.A0N(REG2[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U325 (
	.Y(n210),
	.B1(n159),
	.B0(n366),
	.A1N(n159),
	.A0N(REG3[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U326 (
	.Y(n211),
	.B1(n159),
	.B0(n367),
	.A1N(n159),
	.A0N(REG3[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U327 (
	.Y(n212),
	.B1(n159),
	.B0(n368),
	.A1N(n159),
	.A0N(REG3[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U328 (
	.Y(n213),
	.B1(n159),
	.B0(n369),
	.A1N(n159),
	.A0N(REG3[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U329 (
	.Y(n214),
	.B1(n159),
	.B0(n370),
	.A1N(n159),
	.A0N(REG3[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U330 (
	.Y(n216),
	.B1(n159),
	.B0(n372),
	.A1N(n159),
	.A0N(REG3[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U331 (
	.Y(n217),
	.B1(n159),
	.B0(n373),
	.A1N(n159),
	.A0N(REG3[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U332 (
	.Y(n202),
	.B1(n157),
	.B0(n366),
	.A1N(n157),
	.A0N(REG2[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U333 (
	.Y(n209),
	.B1(n157),
	.B0(n373),
	.A1N(n157),
	.A0N(REG2[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U334 (
	.Y(n215),
	.B1(n159),
	.B0(n371),
	.A1N(n159),
	.A0N(REG3[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U335 (
	.Y(n314),
	.S1(n336),
	.S0(n339),
	.D(REG3[2]),
	.C(REG2[2]),
	.B(REG1[2]),
	.A(REG0[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U336 (
	.Y(n318),
	.S1(n336),
	.S0(n339),
	.D(REG3[3]),
	.C(REG2[3]),
	.B(REG1[3]),
	.A(REG0[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U337 (
	.Y(n322),
	.S1(n336),
	.S0(n340),
	.D(REG3[4]),
	.C(REG2[4]),
	.B(REG1[4]),
	.A(REG0[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U338 (
	.Y(n330),
	.S1(n336),
	.S0(n340),
	.D(REG3[6]),
	.C(REG2[6]),
	.B(REG1[6]),
	.A(REG0[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U339 (
	.Y(n334),
	.S1(n336),
	.S0(n340),
	.D(REG3[7]),
	.C(REG2[7]),
	.B(REG1[7]),
	.A(REG0[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U340 (
	.Y(n141),
	.S1(N11),
	.S0(n338),
	.D(REG3[0]),
	.C(REG2[0]),
	.B(REG1[0]),
	.A(REG0[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U341 (
	.Y(n145),
	.S1(N11),
	.S0(n339),
	.D(REG3[1]),
	.C(REG2[1]),
	.B(REG1[1]),
	.A(REG0[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U342 (
	.Y(n326),
	.S1(n336),
	.S0(n340),
	.D(REG3[5]),
	.C(REG2[5]),
	.B(REG1[5]),
	.A(REG0[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U343 (
	.Y(n140),
	.S1(N11),
	.S0(n338),
	.D(\Reg_file[7][0] ),
	.C(\Reg_file[6][0] ),
	.B(\Reg_file[5][0] ),
	.A(\Reg_file[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U344 (
	.Y(n144),
	.S1(N11),
	.S0(n339),
	.D(\Reg_file[7][1] ),
	.C(\Reg_file[6][1] ),
	.B(\Reg_file[5][1] ),
	.A(\Reg_file[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U345 (
	.Y(n148),
	.S1(n336),
	.S0(n339),
	.D(\Reg_file[7][2] ),
	.C(\Reg_file[6][2] ),
	.B(\Reg_file[5][2] ),
	.A(\Reg_file[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U346 (
	.Y(n317),
	.S1(n336),
	.S0(n339),
	.D(\Reg_file[7][3] ),
	.C(\Reg_file[6][3] ),
	.B(\Reg_file[5][3] ),
	.A(\Reg_file[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U347 (
	.Y(n321),
	.S1(n336),
	.S0(n339),
	.D(\Reg_file[7][4] ),
	.C(\Reg_file[6][4] ),
	.B(\Reg_file[5][4] ),
	.A(\Reg_file[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U348 (
	.Y(n325),
	.S1(n336),
	.S0(n340),
	.D(\Reg_file[7][5] ),
	.C(\Reg_file[6][5] ),
	.B(\Reg_file[5][5] ),
	.A(\Reg_file[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U349 (
	.Y(n329),
	.S1(n336),
	.S0(n340),
	.D(\Reg_file[7][6] ),
	.C(\Reg_file[6][6] ),
	.B(\Reg_file[5][6] ),
	.A(\Reg_file[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U350 (
	.Y(n333),
	.S1(n336),
	.S0(n340),
	.D(\Reg_file[7][7] ),
	.C(\Reg_file[6][7] ),
	.B(\Reg_file[5][7] ),
	.A(\Reg_file[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U351 (
	.Y(n178),
	.B1(n150),
	.B0(N42),
	.A1(n149),
	.A0(R_REG_DATA[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U352 (
	.Y(N42),
	.S1(N12),
	.S0(N13),
	.D(n138),
	.C(n140),
	.B(n139),
	.A(n141), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U353 (
	.Y(n139),
	.S1(N11),
	.S0(n338),
	.D(\Reg_file[11][0] ),
	.C(\Reg_file[10][0] ),
	.B(\Reg_file[9][0] ),
	.A(\Reg_file[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U354 (
	.Y(n138),
	.S1(N11),
	.S0(n338),
	.D(\Reg_file[15][0] ),
	.C(\Reg_file[14][0] ),
	.B(\Reg_file[13][0] ),
	.A(\Reg_file[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U355 (
	.Y(n179),
	.B1(n150),
	.B0(N41),
	.A1(n149),
	.A0(R_REG_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U356 (
	.Y(N41),
	.S1(N12),
	.S0(N13),
	.D(n142),
	.C(n144),
	.B(n143),
	.A(n145), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U357 (
	.Y(n143),
	.S1(n336),
	.S0(n338),
	.D(\Reg_file[11][1] ),
	.C(\Reg_file[10][1] ),
	.B(\Reg_file[9][1] ),
	.A(\Reg_file[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U358 (
	.Y(n142),
	.S1(n336),
	.S0(n338),
	.D(\Reg_file[15][1] ),
	.C(\Reg_file[14][1] ),
	.B(\Reg_file[13][1] ),
	.A(\Reg_file[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U359 (
	.Y(n180),
	.B1(n150),
	.B0(N40),
	.A1(n149),
	.A0(R_REG_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U360 (
	.Y(N40),
	.S1(N12),
	.S0(N13),
	.D(n146),
	.C(n148),
	.B(n147),
	.A(n314), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U361 (
	.Y(n147),
	.S1(n336),
	.S0(n339),
	.D(\Reg_file[11][2] ),
	.C(\Reg_file[10][2] ),
	.B(\Reg_file[9][2] ),
	.A(\Reg_file[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U362 (
	.Y(n146),
	.S1(n336),
	.S0(n339),
	.D(\Reg_file[15][2] ),
	.C(\Reg_file[14][2] ),
	.B(\Reg_file[13][2] ),
	.A(\Reg_file[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U363 (
	.Y(n181),
	.B1(n150),
	.B0(N39),
	.A1(n149),
	.A0(R_REG_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U364 (
	.Y(N39),
	.S1(N12),
	.S0(N13),
	.D(n315),
	.C(n317),
	.B(n316),
	.A(n318), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U365 (
	.Y(n316),
	.S1(n336),
	.S0(n339),
	.D(\Reg_file[11][3] ),
	.C(\Reg_file[10][3] ),
	.B(\Reg_file[9][3] ),
	.A(\Reg_file[8][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U366 (
	.Y(n315),
	.S1(n336),
	.S0(n339),
	.D(\Reg_file[15][3] ),
	.C(\Reg_file[14][3] ),
	.B(\Reg_file[13][3] ),
	.A(\Reg_file[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U367 (
	.Y(n182),
	.B1(n150),
	.B0(N38),
	.A1(n149),
	.A0(R_REG_DATA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U368 (
	.Y(N38),
	.S1(N12),
	.S0(N13),
	.D(n319),
	.C(n321),
	.B(n320),
	.A(n322), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U369 (
	.Y(n320),
	.S1(n336),
	.S0(n339),
	.D(\Reg_file[11][4] ),
	.C(\Reg_file[10][4] ),
	.B(\Reg_file[9][4] ),
	.A(\Reg_file[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U370 (
	.Y(n319),
	.S1(n336),
	.S0(n339),
	.D(\Reg_file[15][4] ),
	.C(\Reg_file[14][4] ),
	.B(\Reg_file[13][4] ),
	.A(\Reg_file[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U371 (
	.Y(n183),
	.B1(n150),
	.B0(N37),
	.A1(n149),
	.A0(R_REG_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U372 (
	.Y(N37),
	.S1(N12),
	.S0(N13),
	.D(n323),
	.C(n325),
	.B(n324),
	.A(n326), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U373 (
	.Y(n324),
	.S1(n336),
	.S0(n340),
	.D(\Reg_file[11][5] ),
	.C(\Reg_file[10][5] ),
	.B(\Reg_file[9][5] ),
	.A(\Reg_file[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U374 (
	.Y(n323),
	.S1(n336),
	.S0(n340),
	.D(\Reg_file[15][5] ),
	.C(\Reg_file[14][5] ),
	.B(\Reg_file[13][5] ),
	.A(\Reg_file[12][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U375 (
	.Y(n184),
	.B1(n150),
	.B0(N36),
	.A1(n149),
	.A0(R_REG_DATA[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U376 (
	.Y(N36),
	.S1(N12),
	.S0(N13),
	.D(n327),
	.C(n329),
	.B(n328),
	.A(n330), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U377 (
	.Y(n328),
	.S1(n336),
	.S0(n340),
	.D(\Reg_file[11][6] ),
	.C(\Reg_file[10][6] ),
	.B(\Reg_file[9][6] ),
	.A(\Reg_file[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U378 (
	.Y(n327),
	.S1(n336),
	.S0(n340),
	.D(\Reg_file[15][6] ),
	.C(\Reg_file[14][6] ),
	.B(\Reg_file[13][6] ),
	.A(\Reg_file[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U379 (
	.Y(n185),
	.B1(n150),
	.B0(N35),
	.A1(n149),
	.A0(R_REG_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U380 (
	.Y(N35),
	.S1(N12),
	.S0(N13),
	.D(n331),
	.C(n333),
	.B(n332),
	.A(n334), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U381 (
	.Y(n332),
	.S1(n336),
	.S0(n340),
	.D(\Reg_file[11][7] ),
	.C(\Reg_file[10][7] ),
	.B(\Reg_file[9][7] ),
	.A(\Reg_file[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U382 (
	.Y(n331),
	.S1(n336),
	.S0(n340),
	.D(\Reg_file[15][7] ),
	.C(\Reg_file[14][7] ),
	.B(\Reg_file[13][7] ),
	.A(\Reg_file[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U383 (
	.Y(n341),
	.A(N10), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U384 (
	.Y(n342),
	.A(N11), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_RTL_DATA_WIDTH8_test_1 (
	ALU_CLK, 
	RST_SYNC_2, 
	ALU_EN, 
	REG0, 
	REG1, 
	ALU_FUNC, 
	ALU_OUT, 
	ALU_OUT_VALID, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input ALU_CLK;
   input RST_SYNC_2;
   input ALU_EN;
   input [7:0] REG0;
   input [7:0] REG1;
   input [3:0] ALU_FUNC;
   output [15:0] ALU_OUT;
   output ALU_OUT_VALID;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN17_SI;
   wire FE_PHN16_SE;
   wire FE_PHN15_SE;
   wire FE_PHN14_SE;
   wire FE_PHN13_SE;
   wire FE_PHN12_SE;
   wire FE_PHN11_SE;
   wire FE_PHN10_SE;
   wire FE_PHN9_SE;
   wire FE_PHN8_SE;
   wire FE_PHN7_SE;
   wire FE_PHN6_SE;
   wire FE_PHN5_SE;
   wire FE_PHN4_SE;
   wire FE_PHN3_SE;
   wire FE_PHN2_SE;
   wire FE_PHN1_SE;
   wire FE_PHN0_SE;
   wire FE_OFN10_n52;
   wire N90;
   wire N91;
   wire N92;
   wire N93;
   wire N94;
   wire N95;
   wire N96;
   wire N97;
   wire N98;
   wire N99;
   wire N100;
   wire N101;
   wire N102;
   wire N103;
   wire N104;
   wire N105;
   wire N106;
   wire N107;
   wire N108;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N113;
   wire N114;
   wire N115;
   wire N116;
   wire N117;
   wire N118;
   wire N119;
   wire N120;
   wire N121;
   wire N122;
   wire N123;
   wire N124;
   wire N125;
   wire N126;
   wire N127;
   wire N128;
   wire N129;
   wire N130;
   wire N131;
   wire N156;
   wire N157;
   wire N158;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire [15:0] ALU_INT;

   // Module instantiations
   DLY1X1M FE_PHC17_SI (
	.Y(FE_PHN17_SI),
	.A(test_si), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M FE_PHC16_SE (
	.Y(FE_PHN16_SE),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M FE_PHC15_SE (
	.Y(FE_PHN15_SE),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M FE_PHC14_SE (
	.Y(FE_PHN14_SE),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M FE_PHC13_SE (
	.Y(FE_PHN13_SE),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M FE_PHC12_SE (
	.Y(FE_PHN12_SE),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M FE_PHC11_SE (
	.Y(FE_PHN11_SE),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M FE_PHC10_SE (
	.Y(FE_PHN10_SE),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M FE_PHC9_SE (
	.Y(FE_PHN9_SE),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M FE_PHC8_SE (
	.Y(FE_PHN8_SE),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M FE_PHC7_SE (
	.Y(FE_PHN7_SE),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M FE_PHC6_SE (
	.Y(FE_PHN6_SE),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M FE_PHC5_SE (
	.Y(FE_PHN5_SE),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M FE_PHC4_SE (
	.Y(FE_PHN4_SE),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X1M FE_PHC3_SE (
	.Y(FE_PHN3_SE),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M FE_PHC2_SE (
	.Y(FE_PHN2_SE),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M FE_PHC1_SE (
	.Y(FE_PHN1_SE),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M FE_PHC0_SE (
	.Y(FE_PHN0_SE),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M FE_OFC10_n52 (
	.Y(FE_OFN10_n52),
	.A(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[15]  (
	.SI(ALU_OUT[14]),
	.SE(FE_PHN16_SE),
	.RN(RST_SYNC_2),
	.Q(ALU_OUT[15]),
	.D(ALU_INT[15]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[14]  (
	.SI(ALU_OUT[13]),
	.SE(FE_PHN5_SE),
	.RN(RST_SYNC_2),
	.Q(ALU_OUT[14]),
	.D(ALU_INT[14]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[13]  (
	.SI(ALU_OUT[12]),
	.SE(FE_PHN6_SE),
	.RN(RST_SYNC_2),
	.Q(ALU_OUT[13]),
	.D(ALU_INT[13]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[12]  (
	.SI(ALU_OUT[11]),
	.SE(FE_PHN4_SE),
	.RN(RST_SYNC_2),
	.Q(ALU_OUT[12]),
	.D(ALU_INT[12]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[11]  (
	.SI(ALU_OUT[10]),
	.SE(FE_PHN2_SE),
	.RN(RST_SYNC_2),
	.Q(ALU_OUT[11]),
	.D(ALU_INT[11]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[10]  (
	.SI(ALU_OUT[9]),
	.SE(FE_PHN1_SE),
	.RN(RST_SYNC_2),
	.Q(ALU_OUT[10]),
	.D(ALU_INT[10]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[9]  (
	.SI(ALU_OUT[8]),
	.SE(FE_PHN3_SE),
	.RN(RST_SYNC_2),
	.Q(ALU_OUT[9]),
	.D(ALU_INT[9]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[8]  (
	.SI(ALU_OUT[7]),
	.SE(FE_PHN12_SE),
	.RN(RST_SYNC_2),
	.Q(ALU_OUT[8]),
	.D(ALU_INT[8]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[7]  (
	.SI(ALU_OUT[6]),
	.SE(FE_PHN11_SE),
	.RN(RST_SYNC_2),
	.Q(ALU_OUT[7]),
	.D(ALU_INT[7]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[6]  (
	.SI(ALU_OUT[5]),
	.SE(FE_PHN14_SE),
	.RN(RST_SYNC_2),
	.Q(ALU_OUT[6]),
	.D(ALU_INT[6]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[5]  (
	.SI(ALU_OUT[4]),
	.SE(FE_PHN13_SE),
	.RN(RST_SYNC_2),
	.Q(ALU_OUT[5]),
	.D(ALU_INT[5]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[4]  (
	.SI(ALU_OUT[3]),
	.SE(FE_PHN10_SE),
	.RN(RST_SYNC_2),
	.Q(ALU_OUT[4]),
	.D(ALU_INT[4]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[3]  (
	.SI(ALU_OUT[2]),
	.SE(FE_PHN9_SE),
	.RN(RST_SYNC_2),
	.Q(ALU_OUT[3]),
	.D(ALU_INT[3]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[2]  (
	.SI(ALU_OUT[1]),
	.SE(FE_PHN8_SE),
	.RN(RST_SYNC_2),
	.Q(ALU_OUT[2]),
	.D(ALU_INT[2]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[1]  (
	.SI(ALU_OUT[0]),
	.SE(FE_PHN7_SE),
	.RN(RST_SYNC_2),
	.Q(ALU_OUT[1]),
	.D(ALU_INT[1]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[0]  (
	.SI(ALU_OUT_VALID),
	.SE(FE_PHN15_SE),
	.RN(RST_SYNC_2),
	.Q(ALU_OUT[0]),
	.D(ALU_INT[0]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M ALU_OUT_VALID_reg (
	.SI(FE_PHN17_SI),
	.SE(FE_PHN0_SE),
	.RN(RST_SYNC_2),
	.Q(ALU_OUT_VALID),
	.D(ALU_EN),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U23 (
	.Y(n64),
	.B0(n118),
	.A1N(n122),
	.A0N(n157), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U24 (
	.Y(n65),
	.B0(n118),
	.A1N(n116),
	.A0N(n117), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U25 (
	.Y(n54),
	.B(n154),
	.AN(n123), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U26 (
	.Y(n59),
	.B(n122),
	.A(n116), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U27 (
	.Y(n48),
	.B(n152),
	.AN(FE_OFN10_n52), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U28 (
	.Y(n67),
	.B(n122),
	.A(n123), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U30 (
	.Y(n58),
	.B(n154),
	.A(n124), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U31 (
	.Y(n154),
	.A(n117), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U32 (
	.Y(n155),
	.A(n108), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U33 (
	.Y(ALU_INT[9]),
	.B0(n49),
	.A1N(n48),
	.A0N(N117), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U34 (
	.Y(ALU_INT[10]),
	.B0(n49),
	.A1N(n48),
	.A0N(N118), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U35 (
	.Y(ALU_INT[11]),
	.B0(n49),
	.A1N(n48),
	.A0N(N119), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U36 (
	.Y(ALU_INT[12]),
	.B0(n49),
	.A1N(n48),
	.A0N(N120), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U37 (
	.Y(ALU_INT[13]),
	.B0(n49),
	.A1N(n48),
	.A0N(N121), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U38 (
	.Y(ALU_INT[14]),
	.B0(n49),
	.A1N(n48),
	.A0N(N122), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U39 (
	.Y(ALU_INT[15]),
	.B0(n49),
	.A1N(n48),
	.A0N(N123), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U40 (
	.Y(n157),
	.A(n124), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3BX2M U41 (
	.Y(n66),
	.C(ALU_FUNC[2]),
	.B(n156),
	.AN(n122), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U42 (
	.Y(n52),
	.C(n156),
	.B(ALU_FUNC[2]),
	.A(n154), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U43 (
	.Y(n123),
	.B(ALU_FUNC[1]),
	.A(ALU_FUNC[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U44 (
	.Y(n63),
	.C(ALU_FUNC[3]),
	.B(n153),
	.A(n123), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U45 (
	.Y(n53),
	.C(ALU_FUNC[3]),
	.B(n153),
	.A(n157), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U46 (
	.Y(n124),
	.B(ALU_FUNC[1]),
	.A(ALU_FUNC[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U47 (
	.Y(n153),
	.A(ALU_FUNC[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U48 (
	.Y(n122),
	.B(ALU_FUNC[3]),
	.A(n153), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U49 (
	.Y(n117),
	.B(ALU_FUNC[0]),
	.A(ALU_FUNC[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U50 (
	.Y(n108),
	.C(n116),
	.B(ALU_FUNC[0]),
	.A(ALU_FUNC[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U51 (
	.Y(n156),
	.A(ALU_FUNC[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U52 (
	.Y(n118),
	.C(ALU_FUNC[3]),
	.B(ALU_FUNC[0]),
	.A(n123), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U53 (
	.Y(n49),
	.B(n140),
	.A(ALU_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U54 (
	.Y(n116),
	.B(n156),
	.A(ALU_FUNC[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U55 (
	.Y(n107),
	.D(n153),
	.C(ALU_FUNC[3]),
	.B(n116),
	.A(N158), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U56 (
	.Y(n152),
	.A(ALU_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U57 (
	.Y(n71),
	.C1(n146),
	.C0(n53),
	.B1(n73),
	.B0(REG1[6]),
	.A1(n139),
	.A0(n72), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U58 (
	.Y(n73),
	.C0(n58),
	.B1(n145),
	.B0(n64),
	.A1(n63),
	.A0(REG0[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U59 (
	.Y(n72),
	.C0(n59),
	.B1(n65),
	.B0(REG0[6]),
	.A1(n145),
	.A0(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U60 (
	.Y(n137),
	.A(n42), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U61 (
	.Y(ALU_INT[2]),
	.B0(n152),
	.A2(n94),
	.A1(n93),
	.A0(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U62 (
	.Y(n92),
	.B1(n54),
	.B0(N92),
	.A1(n67),
	.A0(N101), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U63 (
	.Y(n94),
	.C0(n95),
	.B1(n149),
	.B0(n58),
	.A1(n155),
	.A0(REG0[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U64 (
	.Y(n93),
	.C1(n66),
	.C0(N126),
	.B1(n59),
	.B0(REG0[2]),
	.A1(FE_OFN10_n52),
	.A0(N110), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U65 (
	.Y(ALU_INT[3]),
	.B0(n152),
	.A2(n88),
	.A1(n87),
	.A0(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U66 (
	.Y(n86),
	.B1(n54),
	.B0(N93),
	.A1(n67),
	.A0(N102), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U67 (
	.Y(n88),
	.C0(n89),
	.B1(n148),
	.B0(n58),
	.A1(n155),
	.A0(REG0[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U68 (
	.Y(n87),
	.C1(n66),
	.C0(N127),
	.B1(n59),
	.B0(REG0[3]),
	.A1(FE_OFN10_n52),
	.A0(N111), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U69 (
	.Y(ALU_INT[4]),
	.B0(n152),
	.A2(n82),
	.A1(n81),
	.A0(n80), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U70 (
	.Y(n80),
	.B1(n54),
	.B0(N94),
	.A1(n67),
	.A0(N103), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U71 (
	.Y(n82),
	.C0(n83),
	.B1(n147),
	.B0(n58),
	.A1(REG0[5]),
	.A0(n155), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U72 (
	.Y(n81),
	.C1(n66),
	.C0(N128),
	.B1(n59),
	.B0(REG0[4]),
	.A1(FE_OFN10_n52),
	.A0(N112), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U73 (
	.Y(ALU_INT[5]),
	.B0(n152),
	.A2(n76),
	.A1(n75),
	.A0(n74), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U74 (
	.Y(n74),
	.B1(n54),
	.B0(N95),
	.A1(n67),
	.A0(N104), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U75 (
	.Y(n76),
	.C0(n77),
	.B1(n146),
	.B0(n58),
	.A1(REG0[6]),
	.A0(n155), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U76 (
	.Y(n75),
	.C1(n66),
	.C0(N129),
	.B1(n59),
	.B0(REG0[5]),
	.A1(FE_OFN10_n52),
	.A0(N113), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U77 (
	.Y(ALU_INT[6]),
	.B0(n152),
	.A2(n70),
	.A1(n69),
	.A0(n68), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U78 (
	.Y(n68),
	.B1(n54),
	.B0(N96),
	.A1(n67),
	.A0(N105), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U79 (
	.Y(n70),
	.C0(n71),
	.B1(n145),
	.B0(n58),
	.A1(REG0[7]),
	.A0(n155), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U80 (
	.Y(n69),
	.C1(n66),
	.C0(N130),
	.B1(REG0[6]),
	.B0(n59),
	.A1(FE_OFN10_n52),
	.A0(N114), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U81 (
	.Y(ALU_INT[7]),
	.B0(n152),
	.A2(n57),
	.A1(n56),
	.A0(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U82 (
	.Y(n56),
	.B1(FE_OFN10_n52),
	.B0(N115),
	.A1(n66),
	.A0(N131), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U83 (
	.Y(n55),
	.B1(n54),
	.B0(N97),
	.A1(n67),
	.A0(N106), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U84 (
	.Y(n57),
	.C0(n60),
	.B1(REG0[7]),
	.B0(n59),
	.A1(n144),
	.A0(n58), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U85 (
	.Y(ALU_INT[0]),
	.B0(n152),
	.A2(n112),
	.A1(n111),
	.A0(n110), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U86 (
	.Y(n110),
	.B1(n54),
	.B0(N90),
	.A1(n67),
	.A0(N99), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U87 (
	.Y(n112),
	.C0(n114),
	.B0(n113),
	.A1(n151),
	.A0(n58), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U88 (
	.Y(n111),
	.C1(n66),
	.C0(N124),
	.B1(n59),
	.B0(REG0[0]),
	.A1(FE_OFN10_n52),
	.A0(N108), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U89 (
	.Y(ALU_INT[1]),
	.B0(n152),
	.A2(n100),
	.A1(n99),
	.A0(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U90 (
	.Y(n100),
	.C0(n102),
	.B0(n101),
	.A1(n155),
	.A0(REG0[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U91 (
	.Y(n99),
	.C1(n59),
	.C0(REG0[1]),
	.B1(n150),
	.B0(n58),
	.A1(n66),
	.A0(N125), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U92 (
	.Y(n98),
	.C1(n67),
	.C0(N100),
	.B1(FE_OFN10_n52),
	.B0(N109),
	.A1(n54),
	.A0(N91), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U93 (
	.Y(n140),
	.A(n109), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U94 (
	.Y(n109),
	.C0(n64),
	.B0(n58),
	.A1(n67),
	.A0(N107), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U95 (
	.Y(ALU_INT[8]),
	.B0(n152),
	.A1(n51),
	.A0(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U96 (
	.Y(n50),
	.B0(n140),
	.A1(n54),
	.A0(N98), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB2XLM U97 (
	.Y(n51),
	.B1(FE_OFN10_n52),
	.B0(N116),
	.A1N(n53),
	.A0N(n144), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U98 (
	.Y(N157),
	.A(n133), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U99 (
	.Y(n139),
	.A(REG1[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U101 (
	.Y(n150),
	.A(REG0[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U102 (
	.Y(n151),
	.A(REG0[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U103 (
	.Y(n145),
	.A(REG0[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U104 (
	.Y(n144),
	.A(REG0[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U105 (
	.Y(n148),
	.A(REG0[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U106 (
	.Y(n149),
	.A(REG0[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U107 (
	.Y(n146),
	.A(REG0[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U108 (
	.Y(n147),
	.A(REG0[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U109 (
	.Y(n95),
	.C1(n150),
	.C0(n53),
	.B1(n97),
	.B0(REG1[2]),
	.A1(n136),
	.A0(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U110 (
	.Y(n97),
	.C0(n58),
	.B1(n149),
	.B0(n64),
	.A1(n63),
	.A0(REG0[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U111 (
	.Y(n96),
	.C0(n59),
	.B1(n65),
	.B0(REG0[2]),
	.A1(n149),
	.A0(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U112 (
	.Y(n89),
	.C1(n149),
	.C0(n53),
	.B1(n91),
	.B0(REG1[3]),
	.A1(n138),
	.A0(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U113 (
	.Y(n91),
	.C0(n58),
	.B1(n148),
	.B0(n64),
	.A1(n63),
	.A0(REG0[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U114 (
	.Y(n90),
	.C0(n59),
	.B1(n65),
	.B0(REG0[3]),
	.A1(n148),
	.A0(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U115 (
	.Y(n83),
	.C1(n148),
	.C0(n53),
	.B1(n85),
	.B0(REG1[4]),
	.A1(n143),
	.A0(n84), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U116 (
	.Y(n143),
	.A(REG1[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U117 (
	.Y(n85),
	.C0(n58),
	.B1(n147),
	.B0(n64),
	.A1(n63),
	.A0(REG0[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U118 (
	.Y(n84),
	.C0(n59),
	.B1(n65),
	.B0(REG0[4]),
	.A1(n147),
	.A0(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U119 (
	.Y(n77),
	.C1(n147),
	.C0(n53),
	.B1(n79),
	.B0(REG1[5]),
	.A1(n142),
	.A0(n78), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U120 (
	.Y(n142),
	.A(REG1[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U121 (
	.Y(n79),
	.C0(n58),
	.B1(n146),
	.B0(n64),
	.A1(n63),
	.A0(REG0[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U122 (
	.Y(n78),
	.C0(n59),
	.B1(n65),
	.B0(REG0[5]),
	.A1(n146),
	.A0(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U123 (
	.Y(n60),
	.C1(n145),
	.C0(n53),
	.B1(n62),
	.B0(REG1[7]),
	.A1(n141),
	.A0(n61), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U124 (
	.Y(n141),
	.A(REG1[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U125 (
	.Y(n62),
	.C0(n58),
	.B1(n144),
	.B0(n64),
	.A1(REG0[7]),
	.A0(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U126 (
	.Y(n61),
	.C0(n59),
	.B1(n65),
	.B0(REG0[7]),
	.A1(n144),
	.A0(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U127 (
	.Y(n135),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U128 (
	.Y(n114),
	.B1(n150),
	.B0(n108),
	.A1N(REG1[0]),
	.A0(n115), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U129 (
	.Y(n115),
	.C0(n59),
	.B1(n65),
	.B0(REG0[0]),
	.A1(n151),
	.A0(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U130 (
	.Y(n102),
	.B1(n151),
	.B0(n53),
	.A1N(REG1[1]),
	.A0(n103), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U131 (
	.Y(n103),
	.C0(n59),
	.B1(n65),
	.B0(REG0[1]),
	.A1(n150),
	.A0(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U132 (
	.Y(n113),
	.B0(n120),
	.A1(n119),
	.A0(REG1[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U133 (
	.Y(n120),
	.B0(n107),
	.A2(n121),
	.A1(ALU_FUNC[3]),
	.A0(N156), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U134 (
	.Y(n119),
	.C0(n58),
	.B1(n151),
	.B0(n64),
	.A1(n63),
	.A0(REG0[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U135 (
	.Y(n121),
	.C(ALU_FUNC[0]),
	.B(ALU_FUNC[2]),
	.A(n156), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U136 (
	.Y(n101),
	.B0(n105),
	.A1(n104),
	.A0(REG1[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U137 (
	.Y(n105),
	.B0(n107),
	.A2(n106),
	.A1(ALU_FUNC[3]),
	.A0(N157), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U138 (
	.Y(n104),
	.C0(n58),
	.B1(n150),
	.B0(n64),
	.A1(n63),
	.A0(REG0[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U139 (
	.Y(n106),
	.C(n156),
	.B(ALU_FUNC[2]),
	.A(n153), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U148 (
	.Y(n134),
	.A(REG1[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U149 (
	.Y(n136),
	.A(REG1[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U150 (
	.Y(n138),
	.A(REG1[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U151 (
	.Y(n130),
	.B(REG1[7]),
	.A(n144), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U152 (
	.Y(n46),
	.B(REG0[4]),
	.AN(REG1[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U153 (
	.Y(n35),
	.B(REG1[4]),
	.AN(REG0[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U154 (
	.Y(n125),
	.B(n35),
	.A(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U155 (
	.Y(n43),
	.B(REG0[3]),
	.A(n138), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U156 (
	.Y(n34),
	.B(REG0[2]),
	.A(n136), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U157 (
	.Y(n31),
	.B(REG0[0]),
	.A(n134), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U158 (
	.Y(n45),
	.B(n136),
	.A(REG0[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U159 (
	.Y(n40),
	.B(n45),
	.AN(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X1M U160 (
	.Y(n32),
	.B0(REG1[1]),
	.A1(n150),
	.A0(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X1M U161 (
	.Y(n33),
	.C0(n32),
	.B0(n40),
	.A1(n135),
	.A0(REG0[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U162 (
	.Y(n44),
	.B(n138),
	.A(REG0[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U163 (
	.Y(n36),
	.B0(n44),
	.A2(n33),
	.A1(n34),
	.A0(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U164 (
	.Y(n128),
	.B(REG1[5]),
	.AN(REG0[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X1M U165 (
	.Y(n37),
	.C0(n128),
	.B0(n35),
	.A1(n36),
	.A0(n125), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U166 (
	.Y(n47),
	.B(REG0[5]),
	.AN(REG1[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U167 (
	.Y(n127),
	.B(REG1[6]),
	.A(REG0[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U168 (
	.Y(n38),
	.B1(n145),
	.B0(REG1[6]),
	.A2(n127),
	.A1(n47),
	.A0(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U169 (
	.Y(n131),
	.B(n144),
	.A(REG1[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U170 (
	.Y(N158),
	.B0(n131),
	.A1(n38),
	.A0(n130), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U171 (
	.Y(n41),
	.B(n134),
	.A(REG0[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U172 (
	.Y(n39),
	.B0(REG1[1]),
	.A1(n150),
	.A0(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X1M U173 (
	.Y(n42),
	.C0(n39),
	.B0(n40),
	.A1(n150),
	.A0(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X1M U174 (
	.Y(n126),
	.B0(n43),
	.A2(n44),
	.A1(n45),
	.A0(n137), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X1M U175 (
	.Y(n129),
	.C0(n46),
	.B0(n47),
	.A1N(n126),
	.A0(n125), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U176 (
	.Y(n132),
	.B1(n139),
	.B0(REG0[6]),
	.A2(n127),
	.A1(n128),
	.A0(n129), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X1M U177 (
	.Y(n133),
	.B0(n130),
	.A1N(n132),
	.A0(n131), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U178 (
	.Y(N156),
	.B(N157),
	.A(N158), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_RTL_DATA_WIDTH8_DW_div_uns_0 div_22 (
	.a({ REG0[7],
		REG0[6],
		REG0[5],
		REG0[4],
		REG0[3],
		REG0[2],
		REG0[1],
		REG0[0] }),
	.b({ REG1[7],
		REG1[6],
		REG1[5],
		REG1[4],
		REG1[3],
		REG1[2],
		REG1[1],
		REG1[0] }),
	.quotient({ N131,
		N130,
		N129,
		N128,
		N127,
		N126,
		N125,
		N124 }), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_RTL_DATA_WIDTH8_DW01_sub_0 sub_20 (
	.A({ 1'b0,
		REG0[7],
		REG0[6],
		REG0[5],
		REG0[4],
		REG0[3],
		REG0[2],
		REG0[1],
		REG0[0] }),
	.B({ 1'b0,
		REG1[7],
		REG1[6],
		REG1[5],
		REG1[4],
		REG1[3],
		REG1[2],
		REG1[1],
		REG1[0] }),
	.CI(1'b0),
	.DIFF({ N107,
		N106,
		N105,
		N104,
		N103,
		N102,
		N101,
		N100,
		N99 }), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_RTL_DATA_WIDTH8_DW01_add_0 add_19 (
	.A({ 1'b0,
		REG0[7],
		REG0[6],
		REG0[5],
		REG0[4],
		REG0[3],
		REG0[2],
		REG0[1],
		REG0[0] }),
	.B({ 1'b0,
		REG1[7],
		REG1[6],
		REG1[5],
		REG1[4],
		REG1[3],
		REG1[2],
		REG1[1],
		REG1[0] }),
	.CI(1'b0),
	.SUM({ N98,
		N97,
		N96,
		N95,
		N94,
		N93,
		N92,
		N91,
		N90 }), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_RTL_DATA_WIDTH8_DW02_mult_0 mult_21 (
	.A({ REG0[7],
		REG0[6],
		REG0[5],
		REG0[4],
		REG0[3],
		REG0[2],
		REG0[1],
		REG0[0] }),
	.B({ REG1[7],
		REG1[6],
		REG1[5],
		REG1[4],
		REG1[3],
		REG1[2],
		REG1[1],
		REG1[0] }),
	.TC(1'b0),
	.PRODUCT({ N123,
		N122,
		N121,
		N120,
		N119,
		N118,
		N117,
		N116,
		N115,
		N114,
		N113,
		N112,
		N111,
		N110,
		N109,
		N108 }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_RTL_DATA_WIDTH8_DW_div_uns_0 (
	a, 
	b, 
	quotient, 
	remainder, 
	divide_by_0, 
	VDD, 
	VSS);
   input [7:0] a;
   input [7:0] b;
   output [7:0] quotient;
   output [7:0] remainder;
   output divide_by_0;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \u_div/SumTmp[1][0] ;
   wire \u_div/SumTmp[1][1] ;
   wire \u_div/SumTmp[1][2] ;
   wire \u_div/SumTmp[1][3] ;
   wire \u_div/SumTmp[1][4] ;
   wire \u_div/SumTmp[1][5] ;
   wire \u_div/SumTmp[1][6] ;
   wire \u_div/SumTmp[2][0] ;
   wire \u_div/SumTmp[2][1] ;
   wire \u_div/SumTmp[2][2] ;
   wire \u_div/SumTmp[2][3] ;
   wire \u_div/SumTmp[2][4] ;
   wire \u_div/SumTmp[2][5] ;
   wire \u_div/SumTmp[3][0] ;
   wire \u_div/SumTmp[3][1] ;
   wire \u_div/SumTmp[3][2] ;
   wire \u_div/SumTmp[3][3] ;
   wire \u_div/SumTmp[3][4] ;
   wire \u_div/SumTmp[4][0] ;
   wire \u_div/SumTmp[4][1] ;
   wire \u_div/SumTmp[4][2] ;
   wire \u_div/SumTmp[4][3] ;
   wire \u_div/SumTmp[5][0] ;
   wire \u_div/SumTmp[5][1] ;
   wire \u_div/SumTmp[5][2] ;
   wire \u_div/SumTmp[6][0] ;
   wire \u_div/SumTmp[6][1] ;
   wire \u_div/SumTmp[7][0] ;
   wire \u_div/CryTmp[0][1] ;
   wire \u_div/CryTmp[0][2] ;
   wire \u_div/CryTmp[0][3] ;
   wire \u_div/CryTmp[0][4] ;
   wire \u_div/CryTmp[0][5] ;
   wire \u_div/CryTmp[0][6] ;
   wire \u_div/CryTmp[0][7] ;
   wire \u_div/CryTmp[1][1] ;
   wire \u_div/CryTmp[1][2] ;
   wire \u_div/CryTmp[1][3] ;
   wire \u_div/CryTmp[1][4] ;
   wire \u_div/CryTmp[1][5] ;
   wire \u_div/CryTmp[1][6] ;
   wire \u_div/CryTmp[1][7] ;
   wire \u_div/CryTmp[2][1] ;
   wire \u_div/CryTmp[2][2] ;
   wire \u_div/CryTmp[2][3] ;
   wire \u_div/CryTmp[2][4] ;
   wire \u_div/CryTmp[2][5] ;
   wire \u_div/CryTmp[2][6] ;
   wire \u_div/CryTmp[3][1] ;
   wire \u_div/CryTmp[3][2] ;
   wire \u_div/CryTmp[3][3] ;
   wire \u_div/CryTmp[3][4] ;
   wire \u_div/CryTmp[3][5] ;
   wire \u_div/CryTmp[4][1] ;
   wire \u_div/CryTmp[4][2] ;
   wire \u_div/CryTmp[4][3] ;
   wire \u_div/CryTmp[4][4] ;
   wire \u_div/CryTmp[5][1] ;
   wire \u_div/CryTmp[5][2] ;
   wire \u_div/CryTmp[5][3] ;
   wire \u_div/CryTmp[6][1] ;
   wire \u_div/CryTmp[6][2] ;
   wire \u_div/CryTmp[7][1] ;
   wire \u_div/PartRem[1][1] ;
   wire \u_div/PartRem[1][2] ;
   wire \u_div/PartRem[1][3] ;
   wire \u_div/PartRem[1][4] ;
   wire \u_div/PartRem[1][5] ;
   wire \u_div/PartRem[1][6] ;
   wire \u_div/PartRem[1][7] ;
   wire \u_div/PartRem[2][1] ;
   wire \u_div/PartRem[2][2] ;
   wire \u_div/PartRem[2][3] ;
   wire \u_div/PartRem[2][4] ;
   wire \u_div/PartRem[2][5] ;
   wire \u_div/PartRem[2][6] ;
   wire \u_div/PartRem[3][1] ;
   wire \u_div/PartRem[3][2] ;
   wire \u_div/PartRem[3][3] ;
   wire \u_div/PartRem[3][4] ;
   wire \u_div/PartRem[3][5] ;
   wire \u_div/PartRem[4][1] ;
   wire \u_div/PartRem[4][2] ;
   wire \u_div/PartRem[4][3] ;
   wire \u_div/PartRem[4][4] ;
   wire \u_div/PartRem[5][1] ;
   wire \u_div/PartRem[5][2] ;
   wire \u_div/PartRem[5][3] ;
   wire \u_div/PartRem[6][1] ;
   wire \u_div/PartRem[6][2] ;
   wire \u_div/PartRem[7][1] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;

   // Module instantiations
   ADDFX2M \u_div/u_fa_PartRem_0_2_5  (
	.S(\u_div/SumTmp[2][5] ),
	.CO(\u_div/CryTmp[2][6] ),
	.CI(\u_div/CryTmp[2][5] ),
	.B(n13),
	.A(\u_div/PartRem[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_4_3  (
	.S(\u_div/SumTmp[4][3] ),
	.CO(\u_div/CryTmp[4][4] ),
	.CI(\u_div/CryTmp[4][3] ),
	.B(n15),
	.A(\u_div/PartRem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_5_2  (
	.S(\u_div/SumTmp[5][2] ),
	.CO(\u_div/CryTmp[5][3] ),
	.CI(\u_div/CryTmp[5][2] ),
	.B(n16),
	.A(\u_div/PartRem[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_6_1  (
	.S(\u_div/SumTmp[6][1] ),
	.CO(\u_div/CryTmp[6][2] ),
	.CI(\u_div/CryTmp[6][1] ),
	.B(n17),
	.A(\u_div/PartRem[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_3_4  (
	.S(\u_div/SumTmp[3][4] ),
	.CO(\u_div/CryTmp[3][5] ),
	.CI(\u_div/CryTmp[3][4] ),
	.B(n14),
	.A(\u_div/PartRem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_5  (
	.CO(\u_div/CryTmp[0][6] ),
	.CI(\u_div/CryTmp[0][5] ),
	.B(n13),
	.A(\u_div/PartRem[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_6  (
	.CO(\u_div/CryTmp[0][7] ),
	.CI(\u_div/CryTmp[0][6] ),
	.B(n12),
	.A(\u_div/PartRem[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_7  (
	.CO(quotient[0]),
	.CI(\u_div/CryTmp[0][7] ),
	.B(n11),
	.A(\u_div/PartRem[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_1  (
	.CO(\u_div/CryTmp[0][2] ),
	.CI(\u_div/CryTmp[0][1] ),
	.B(n17),
	.A(\u_div/PartRem[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_1  (
	.S(\u_div/SumTmp[1][1] ),
	.CO(\u_div/CryTmp[1][2] ),
	.CI(\u_div/CryTmp[1][1] ),
	.B(n17),
	.A(\u_div/PartRem[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_2_1  (
	.S(\u_div/SumTmp[2][1] ),
	.CO(\u_div/CryTmp[2][2] ),
	.CI(\u_div/CryTmp[2][1] ),
	.B(n17),
	.A(\u_div/PartRem[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_3_1  (
	.S(\u_div/SumTmp[3][1] ),
	.CO(\u_div/CryTmp[3][2] ),
	.CI(\u_div/CryTmp[3][1] ),
	.B(n17),
	.A(\u_div/PartRem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_4_1  (
	.S(\u_div/SumTmp[4][1] ),
	.CO(\u_div/CryTmp[4][2] ),
	.CI(\u_div/CryTmp[4][1] ),
	.B(n17),
	.A(\u_div/PartRem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_5_1  (
	.S(\u_div/SumTmp[5][1] ),
	.CO(\u_div/CryTmp[5][2] ),
	.CI(\u_div/CryTmp[5][1] ),
	.B(n17),
	.A(\u_div/PartRem[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_2  (
	.CO(\u_div/CryTmp[0][3] ),
	.CI(\u_div/CryTmp[0][2] ),
	.B(n16),
	.A(\u_div/PartRem[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_3  (
	.CO(\u_div/CryTmp[0][4] ),
	.CI(\u_div/CryTmp[0][3] ),
	.B(n15),
	.A(\u_div/PartRem[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_4  (
	.CO(\u_div/CryTmp[0][5] ),
	.CI(\u_div/CryTmp[0][4] ),
	.B(n14),
	.A(\u_div/PartRem[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_5  (
	.S(\u_div/SumTmp[1][5] ),
	.CO(\u_div/CryTmp[1][6] ),
	.CI(\u_div/CryTmp[1][5] ),
	.B(n13),
	.A(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_4  (
	.S(\u_div/SumTmp[1][4] ),
	.CO(\u_div/CryTmp[1][5] ),
	.CI(\u_div/CryTmp[1][4] ),
	.B(n14),
	.A(\u_div/PartRem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_3  (
	.S(\u_div/SumTmp[1][3] ),
	.CO(\u_div/CryTmp[1][4] ),
	.CI(\u_div/CryTmp[1][3] ),
	.B(n15),
	.A(\u_div/PartRem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_2_4  (
	.S(\u_div/SumTmp[2][4] ),
	.CO(\u_div/CryTmp[2][5] ),
	.CI(\u_div/CryTmp[2][4] ),
	.B(n14),
	.A(\u_div/PartRem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_2  (
	.S(\u_div/SumTmp[1][2] ),
	.CO(\u_div/CryTmp[1][3] ),
	.CI(\u_div/CryTmp[1][2] ),
	.B(n16),
	.A(\u_div/PartRem[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_2_3  (
	.S(\u_div/SumTmp[2][3] ),
	.CO(\u_div/CryTmp[2][4] ),
	.CI(\u_div/CryTmp[2][3] ),
	.B(n15),
	.A(\u_div/PartRem[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_2_2  (
	.S(\u_div/SumTmp[2][2] ),
	.CO(\u_div/CryTmp[2][3] ),
	.CI(\u_div/CryTmp[2][2] ),
	.B(n16),
	.A(\u_div/PartRem[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_3_3  (
	.S(\u_div/SumTmp[3][3] ),
	.CO(\u_div/CryTmp[3][4] ),
	.CI(\u_div/CryTmp[3][3] ),
	.B(n15),
	.A(\u_div/PartRem[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_3_2  (
	.S(\u_div/SumTmp[3][2] ),
	.CO(\u_div/CryTmp[3][3] ),
	.CI(\u_div/CryTmp[3][2] ),
	.B(n16),
	.A(\u_div/PartRem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_4_2  (
	.S(\u_div/SumTmp[4][2] ),
	.CO(\u_div/CryTmp[4][3] ),
	.CI(\u_div/CryTmp[4][2] ),
	.B(n16),
	.A(\u_div/PartRem[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_6  (
	.S(\u_div/SumTmp[1][6] ),
	.CO(\u_div/CryTmp[1][7] ),
	.CI(\u_div/CryTmp[1][6] ),
	.B(n12),
	.A(\u_div/PartRem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U1 (
	.Y(n18),
	.A(b[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U2 (
	.Y(\u_div/SumTmp[7][0] ),
	.B(a[7]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U3 (
	.Y(\u_div/SumTmp[6][0] ),
	.B(a[6]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U4 (
	.Y(\u_div/SumTmp[5][0] ),
	.B(a[5]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U5 (
	.Y(\u_div/SumTmp[4][0] ),
	.B(a[4]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U6 (
	.Y(\u_div/SumTmp[3][0] ),
	.B(a[3]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U7 (
	.Y(\u_div/SumTmp[2][0] ),
	.B(a[2]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U8 (
	.Y(\u_div/CryTmp[7][1] ),
	.B(a[7]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U9 (
	.Y(\u_div/SumTmp[1][0] ),
	.B(a[1]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U10 (
	.Y(\u_div/CryTmp[5][1] ),
	.B(n3),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U11 (
	.Y(n3),
	.A(a[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(n2),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U13 (
	.Y(\u_div/CryTmp[4][1] ),
	.B(n5),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U14 (
	.Y(n5),
	.A(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U15 (
	.Y(n4),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U16 (
	.Y(\u_div/CryTmp[3][1] ),
	.B(n7),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n7),
	.A(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(n6),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U19 (
	.Y(\u_div/CryTmp[2][1] ),
	.B(n8),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n8),
	.A(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U21 (
	.Y(\u_div/CryTmp[1][1] ),
	.B(n9),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n9),
	.A(a[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U23 (
	.Y(\u_div/CryTmp[0][1] ),
	.B(n10),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U24 (
	.Y(n10),
	.A(a[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U25 (
	.Y(\u_div/CryTmp[6][1] ),
	.B(n1),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U26 (
	.Y(n1),
	.A(a[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U27 (
	.Y(n12),
	.A(b[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U28 (
	.Y(n17),
	.A(b[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U29 (
	.Y(n16),
	.A(b[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U30 (
	.Y(n15),
	.A(b[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U31 (
	.Y(n14),
	.A(b[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U32 (
	.Y(n13),
	.A(b[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U33 (
	.Y(n11),
	.A(b[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U34 (
	.Y(\u_div/PartRem[1][7] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][6] ),
	.A(\u_div/PartRem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U35 (
	.Y(\u_div/PartRem[2][6] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][5] ),
	.A(\u_div/PartRem[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U36 (
	.Y(\u_div/PartRem[3][5] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][4] ),
	.A(\u_div/PartRem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U37 (
	.Y(\u_div/PartRem[4][4] ),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][3] ),
	.A(\u_div/PartRem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U38 (
	.Y(\u_div/PartRem[5][3] ),
	.S0(quotient[5]),
	.B(\u_div/SumTmp[5][2] ),
	.A(\u_div/PartRem[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U39 (
	.Y(\u_div/PartRem[6][2] ),
	.S0(quotient[6]),
	.B(\u_div/SumTmp[6][1] ),
	.A(\u_div/PartRem[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U40 (
	.Y(\u_div/PartRem[7][1] ),
	.S0(quotient[7]),
	.B(\u_div/SumTmp[7][0] ),
	.A(a[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U41 (
	.Y(\u_div/PartRem[1][6] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][5] ),
	.A(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U42 (
	.Y(\u_div/PartRem[2][5] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][4] ),
	.A(\u_div/PartRem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U43 (
	.Y(\u_div/PartRem[3][4] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][3] ),
	.A(\u_div/PartRem[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U44 (
	.Y(\u_div/PartRem[4][3] ),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][2] ),
	.A(\u_div/PartRem[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U45 (
	.Y(\u_div/PartRem[5][2] ),
	.S0(quotient[5]),
	.B(\u_div/SumTmp[5][1] ),
	.A(\u_div/PartRem[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U46 (
	.Y(\u_div/PartRem[6][1] ),
	.S0(quotient[6]),
	.B(\u_div/SumTmp[6][0] ),
	.A(a[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U47 (
	.Y(\u_div/PartRem[1][5] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][4] ),
	.A(\u_div/PartRem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U48 (
	.Y(\u_div/PartRem[2][4] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][3] ),
	.A(\u_div/PartRem[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U49 (
	.Y(\u_div/PartRem[3][3] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][2] ),
	.A(\u_div/PartRem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U50 (
	.Y(\u_div/PartRem[4][2] ),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][1] ),
	.A(\u_div/PartRem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U51 (
	.Y(\u_div/PartRem[5][1] ),
	.S0(quotient[5]),
	.B(\u_div/SumTmp[5][0] ),
	.A(a[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U52 (
	.Y(\u_div/PartRem[1][4] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][3] ),
	.A(\u_div/PartRem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U53 (
	.Y(\u_div/PartRem[2][3] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][2] ),
	.A(\u_div/PartRem[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U54 (
	.Y(\u_div/PartRem[3][2] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][1] ),
	.A(\u_div/PartRem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U55 (
	.Y(\u_div/PartRem[4][1] ),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][0] ),
	.A(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U56 (
	.Y(\u_div/PartRem[1][3] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][2] ),
	.A(\u_div/PartRem[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U57 (
	.Y(\u_div/PartRem[2][2] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][1] ),
	.A(\u_div/PartRem[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U58 (
	.Y(\u_div/PartRem[3][1] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][0] ),
	.A(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U59 (
	.Y(\u_div/PartRem[1][2] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][1] ),
	.A(\u_div/PartRem[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U60 (
	.Y(\u_div/PartRem[2][1] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][0] ),
	.A(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U61 (
	.Y(\u_div/PartRem[1][1] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][0] ),
	.A(a[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X1M U62 (
	.Y(quotient[7]),
	.D(n16),
	.C(n17),
	.B(n19),
	.A(\u_div/CryTmp[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X1M U63 (
	.Y(quotient[6]),
	.C(\u_div/CryTmp[6][2] ),
	.B(n16),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U64 (
	.Y(quotient[5]),
	.B(n19),
	.A(\u_div/CryTmp[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U65 (
	.Y(n19),
	.B(n15),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U66 (
	.Y(quotient[4]),
	.B(n20),
	.A(\u_div/CryTmp[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X1M U67 (
	.Y(n20),
	.C(n13),
	.B(n14),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X1M U68 (
	.Y(quotient[3]),
	.C(\u_div/CryTmp[3][5] ),
	.B(n13),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U69 (
	.Y(quotient[2]),
	.B(n21),
	.A(\u_div/CryTmp[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U70 (
	.Y(n21),
	.B(b[7]),
	.A(b[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U71 (
	.Y(quotient[1]),
	.B(n11),
	.A(\u_div/CryTmp[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_RTL_DATA_WIDTH8_DW01_sub_0 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO, 
	VDD, 
	VSS);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] DIFF;
   output CO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire [9:0] carry;

   // Module instantiations
   ADDFX2M U2_1 (
	.S(DIFF[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(n9),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_5 (
	.S(DIFF[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(n5),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_4 (
	.S(DIFF[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(n6),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_3 (
	.S(DIFF[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(n7),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_2 (
	.S(DIFF[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(n8),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_7 (
	.S(DIFF[7]),
	.CO(carry[8]),
	.CI(carry[7]),
	.B(n3),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_6 (
	.S(DIFF[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(n4),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U1 (
	.Y(DIFF[0]),
	.B(A[0]),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U2 (
	.Y(DIFF[8]),
	.A(carry[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(n4),
	.A(B[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U4 (
	.Y(n10),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(n3),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U6 (
	.Y(n8),
	.A(B[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U7 (
	.Y(n7),
	.A(B[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(n6),
	.A(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U9 (
	.Y(n5),
	.A(B[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U10 (
	.Y(carry[1]),
	.B(n1),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U11 (
	.Y(n9),
	.A(B[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(n1),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_RTL_DATA_WIDTH8_DW01_add_0 (
	A, 
	B, 
	CI, 
	SUM, 
	CO, 
	VDD, 
	VSS);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] SUM;
   output CO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire [8:1] carry;

   // Module instantiations
   ADDFX2M U1_7 (
	.S(SUM[7]),
	.CO(SUM[8]),
	.CI(carry[7]),
	.B(B[7]),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(n1),
	.B(B[1]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U1 (
	.Y(n1),
	.B(A[0]),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U2 (
	.Y(SUM[0]),
	.B(A[0]),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_RTL_DATA_WIDTH8_DW02_mult_0 (
	A, 
	B, 
	TC, 
	PRODUCT, 
	VDD, 
	VSS);
   input [7:0] A;
   input [7:0] B;
   input TC;
   output [15:0] PRODUCT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \ab[7][7] ;
   wire \ab[7][6] ;
   wire \ab[7][5] ;
   wire \ab[7][4] ;
   wire \ab[7][3] ;
   wire \ab[7][2] ;
   wire \ab[7][1] ;
   wire \ab[7][0] ;
   wire \ab[6][7] ;
   wire \ab[6][6] ;
   wire \ab[6][5] ;
   wire \ab[6][4] ;
   wire \ab[6][3] ;
   wire \ab[6][2] ;
   wire \ab[6][1] ;
   wire \ab[6][0] ;
   wire \ab[5][7] ;
   wire \ab[5][6] ;
   wire \ab[5][5] ;
   wire \ab[5][4] ;
   wire \ab[5][3] ;
   wire \ab[5][2] ;
   wire \ab[5][1] ;
   wire \ab[5][0] ;
   wire \ab[4][7] ;
   wire \ab[4][6] ;
   wire \ab[4][5] ;
   wire \ab[4][4] ;
   wire \ab[4][3] ;
   wire \ab[4][2] ;
   wire \ab[4][1] ;
   wire \ab[4][0] ;
   wire \ab[3][7] ;
   wire \ab[3][6] ;
   wire \ab[3][5] ;
   wire \ab[3][4] ;
   wire \ab[3][3] ;
   wire \ab[3][2] ;
   wire \ab[3][1] ;
   wire \ab[3][0] ;
   wire \ab[2][7] ;
   wire \ab[2][6] ;
   wire \ab[2][5] ;
   wire \ab[2][4] ;
   wire \ab[2][3] ;
   wire \ab[2][2] ;
   wire \ab[2][1] ;
   wire \ab[2][0] ;
   wire \ab[1][7] ;
   wire \ab[1][6] ;
   wire \ab[1][5] ;
   wire \ab[1][4] ;
   wire \ab[1][3] ;
   wire \ab[1][2] ;
   wire \ab[1][1] ;
   wire \ab[1][0] ;
   wire \ab[0][7] ;
   wire \ab[0][6] ;
   wire \ab[0][5] ;
   wire \ab[0][4] ;
   wire \ab[0][3] ;
   wire \ab[0][2] ;
   wire \ab[0][1] ;
   wire \CARRYB[7][6] ;
   wire \CARRYB[7][5] ;
   wire \CARRYB[7][4] ;
   wire \CARRYB[7][3] ;
   wire \CARRYB[7][2] ;
   wire \CARRYB[7][1] ;
   wire \CARRYB[7][0] ;
   wire \CARRYB[6][6] ;
   wire \CARRYB[6][5] ;
   wire \CARRYB[6][4] ;
   wire \CARRYB[6][3] ;
   wire \CARRYB[6][2] ;
   wire \CARRYB[6][1] ;
   wire \CARRYB[6][0] ;
   wire \CARRYB[5][6] ;
   wire \CARRYB[5][5] ;
   wire \CARRYB[5][4] ;
   wire \CARRYB[5][3] ;
   wire \CARRYB[5][2] ;
   wire \CARRYB[5][1] ;
   wire \CARRYB[5][0] ;
   wire \CARRYB[4][6] ;
   wire \CARRYB[4][5] ;
   wire \CARRYB[4][4] ;
   wire \CARRYB[4][3] ;
   wire \CARRYB[4][2] ;
   wire \CARRYB[4][1] ;
   wire \CARRYB[4][0] ;
   wire \CARRYB[3][6] ;
   wire \CARRYB[3][5] ;
   wire \CARRYB[3][4] ;
   wire \CARRYB[3][3] ;
   wire \CARRYB[3][2] ;
   wire \CARRYB[3][1] ;
   wire \CARRYB[3][0] ;
   wire \CARRYB[2][6] ;
   wire \CARRYB[2][5] ;
   wire \CARRYB[2][4] ;
   wire \CARRYB[2][3] ;
   wire \CARRYB[2][2] ;
   wire \CARRYB[2][1] ;
   wire \CARRYB[2][0] ;
   wire \SUMB[7][6] ;
   wire \SUMB[7][5] ;
   wire \SUMB[7][4] ;
   wire \SUMB[7][3] ;
   wire \SUMB[7][2] ;
   wire \SUMB[7][1] ;
   wire \SUMB[7][0] ;
   wire \SUMB[6][6] ;
   wire \SUMB[6][5] ;
   wire \SUMB[6][4] ;
   wire \SUMB[6][3] ;
   wire \SUMB[6][2] ;
   wire \SUMB[6][1] ;
   wire \SUMB[5][6] ;
   wire \SUMB[5][5] ;
   wire \SUMB[5][4] ;
   wire \SUMB[5][3] ;
   wire \SUMB[5][2] ;
   wire \SUMB[5][1] ;
   wire \SUMB[4][6] ;
   wire \SUMB[4][5] ;
   wire \SUMB[4][4] ;
   wire \SUMB[4][3] ;
   wire \SUMB[4][2] ;
   wire \SUMB[4][1] ;
   wire \SUMB[3][6] ;
   wire \SUMB[3][5] ;
   wire \SUMB[3][4] ;
   wire \SUMB[3][3] ;
   wire \SUMB[3][2] ;
   wire \SUMB[3][1] ;
   wire \SUMB[2][6] ;
   wire \SUMB[2][5] ;
   wire \SUMB[2][4] ;
   wire \SUMB[2][3] ;
   wire \SUMB[2][2] ;
   wire \SUMB[2][1] ;
   wire \SUMB[1][6] ;
   wire \SUMB[1][5] ;
   wire \SUMB[1][4] ;
   wire \SUMB[1][3] ;
   wire \SUMB[1][2] ;
   wire \SUMB[1][1] ;
   wire \A1[12] ;
   wire \A1[11] ;
   wire \A1[10] ;
   wire \A1[9] ;
   wire \A1[8] ;
   wire \A1[7] ;
   wire \A1[6] ;
   wire \A1[4] ;
   wire \A1[3] ;
   wire \A1[2] ;
   wire \A1[1] ;
   wire \A1[0] ;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;

   // Module instantiations
   ADDFX2M S1_6_0 (
	.S(\A1[4] ),
	.CO(\CARRYB[6][0] ),
	.CI(\SUMB[5][1] ),
	.B(\CARRYB[5][0] ),
	.A(\ab[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_5_0 (
	.S(\A1[3] ),
	.CO(\CARRYB[5][0] ),
	.CI(\SUMB[4][1] ),
	.B(\CARRYB[4][0] ),
	.A(\ab[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_4_0 (
	.S(\A1[2] ),
	.CO(\CARRYB[4][0] ),
	.CI(\SUMB[3][1] ),
	.B(\CARRYB[3][0] ),
	.A(\ab[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_3_0 (
	.S(\A1[1] ),
	.CO(\CARRYB[3][0] ),
	.CI(\SUMB[2][1] ),
	.B(\CARRYB[2][0] ),
	.A(\ab[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_5 (
	.S(\SUMB[6][5] ),
	.CO(\CARRYB[6][5] ),
	.CI(\SUMB[5][6] ),
	.B(\CARRYB[5][5] ),
	.A(\ab[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_4 (
	.S(\SUMB[6][4] ),
	.CO(\CARRYB[6][4] ),
	.CI(\SUMB[5][5] ),
	.B(\CARRYB[5][4] ),
	.A(\ab[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_5 (
	.S(\SUMB[5][5] ),
	.CO(\CARRYB[5][5] ),
	.CI(\SUMB[4][6] ),
	.B(\CARRYB[4][5] ),
	.A(\ab[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_3 (
	.S(\SUMB[6][3] ),
	.CO(\CARRYB[6][3] ),
	.CI(\SUMB[5][4] ),
	.B(\CARRYB[5][3] ),
	.A(\ab[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_4 (
	.S(\SUMB[5][4] ),
	.CO(\CARRYB[5][4] ),
	.CI(\SUMB[4][5] ),
	.B(\CARRYB[4][4] ),
	.A(\ab[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_1 (
	.S(\SUMB[6][1] ),
	.CO(\CARRYB[6][1] ),
	.CI(\SUMB[5][2] ),
	.B(\CARRYB[5][1] ),
	.A(\ab[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_2 (
	.S(\SUMB[6][2] ),
	.CO(\CARRYB[6][2] ),
	.CI(\SUMB[5][3] ),
	.B(\CARRYB[5][2] ),
	.A(\ab[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_5 (
	.S(\SUMB[4][5] ),
	.CO(\CARRYB[4][5] ),
	.CI(\SUMB[3][6] ),
	.B(\CARRYB[3][5] ),
	.A(\ab[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_1 (
	.S(\SUMB[5][1] ),
	.CO(\CARRYB[5][1] ),
	.CI(\SUMB[4][2] ),
	.B(\CARRYB[4][1] ),
	.A(\ab[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_2 (
	.S(\SUMB[5][2] ),
	.CO(\CARRYB[5][2] ),
	.CI(\SUMB[4][3] ),
	.B(\CARRYB[4][2] ),
	.A(\ab[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_3 (
	.S(\SUMB[5][3] ),
	.CO(\CARRYB[5][3] ),
	.CI(\SUMB[4][4] ),
	.B(\CARRYB[4][3] ),
	.A(\ab[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_1 (
	.S(\SUMB[4][1] ),
	.CO(\CARRYB[4][1] ),
	.CI(\SUMB[3][2] ),
	.B(\CARRYB[3][1] ),
	.A(\ab[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_2 (
	.S(\SUMB[4][2] ),
	.CO(\CARRYB[4][2] ),
	.CI(\SUMB[3][3] ),
	.B(\CARRYB[3][2] ),
	.A(\ab[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_3 (
	.S(\SUMB[4][3] ),
	.CO(\CARRYB[4][3] ),
	.CI(\SUMB[3][4] ),
	.B(\CARRYB[3][3] ),
	.A(\ab[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_4 (
	.S(\SUMB[4][4] ),
	.CO(\CARRYB[4][4] ),
	.CI(\SUMB[3][5] ),
	.B(\CARRYB[3][4] ),
	.A(\ab[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_1 (
	.S(\SUMB[3][1] ),
	.CO(\CARRYB[3][1] ),
	.CI(\SUMB[2][2] ),
	.B(\CARRYB[2][1] ),
	.A(\ab[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_2 (
	.S(\SUMB[3][2] ),
	.CO(\CARRYB[3][2] ),
	.CI(\SUMB[2][3] ),
	.B(\CARRYB[2][2] ),
	.A(\ab[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_3 (
	.S(\SUMB[3][3] ),
	.CO(\CARRYB[3][3] ),
	.CI(\SUMB[2][4] ),
	.B(\CARRYB[2][3] ),
	.A(\ab[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_4 (
	.S(\SUMB[3][4] ),
	.CO(\CARRYB[3][4] ),
	.CI(\SUMB[2][5] ),
	.B(\CARRYB[2][4] ),
	.A(\ab[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_5 (
	.S(\SUMB[3][5] ),
	.CO(\CARRYB[3][5] ),
	.CI(\SUMB[2][6] ),
	.B(\CARRYB[2][5] ),
	.A(\ab[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_6_6 (
	.S(\SUMB[6][6] ),
	.CO(\CARRYB[6][6] ),
	.CI(\ab[5][7] ),
	.B(\CARRYB[5][6] ),
	.A(\ab[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_5_6 (
	.S(\SUMB[5][6] ),
	.CO(\CARRYB[5][6] ),
	.CI(\ab[4][7] ),
	.B(\CARRYB[4][6] ),
	.A(\ab[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_4_6 (
	.S(\SUMB[4][6] ),
	.CO(\CARRYB[4][6] ),
	.CI(\ab[3][7] ),
	.B(\CARRYB[3][6] ),
	.A(\ab[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_3_6 (
	.S(\SUMB[3][6] ),
	.CO(\CARRYB[3][6] ),
	.CI(\ab[2][7] ),
	.B(\CARRYB[2][6] ),
	.A(\ab[3][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_2_6 (
	.S(\SUMB[2][6] ),
	.CO(\CARRYB[2][6] ),
	.CI(\ab[1][7] ),
	.B(n8),
	.A(\ab[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_2_0 (
	.S(\A1[0] ),
	.CO(\CARRYB[2][0] ),
	.CI(\SUMB[1][1] ),
	.B(n9),
	.A(\ab[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_1 (
	.S(\SUMB[2][1] ),
	.CO(\CARRYB[2][1] ),
	.CI(\SUMB[1][2] ),
	.B(n7),
	.A(\ab[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_2 (
	.S(\SUMB[2][2] ),
	.CO(\CARRYB[2][2] ),
	.CI(\SUMB[1][3] ),
	.B(n6),
	.A(\ab[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_3 (
	.S(\SUMB[2][3] ),
	.CO(\CARRYB[2][3] ),
	.CI(\SUMB[1][4] ),
	.B(n5),
	.A(\ab[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_4 (
	.S(\SUMB[2][4] ),
	.CO(\CARRYB[2][4] ),
	.CI(\SUMB[1][5] ),
	.B(n4),
	.A(\ab[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_5 (
	.S(\SUMB[2][5] ),
	.CO(\CARRYB[2][5] ),
	.CI(\SUMB[1][6] ),
	.B(n3),
	.A(\ab[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_0 (
	.S(\SUMB[7][0] ),
	.CO(\CARRYB[7][0] ),
	.CI(\SUMB[6][1] ),
	.B(\CARRYB[6][0] ),
	.A(\ab[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S5_6 (
	.S(\SUMB[7][6] ),
	.CO(\CARRYB[7][6] ),
	.CI(\ab[6][7] ),
	.B(\CARRYB[6][6] ),
	.A(\ab[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_5 (
	.S(\SUMB[7][5] ),
	.CO(\CARRYB[7][5] ),
	.CI(\SUMB[6][6] ),
	.B(\CARRYB[6][5] ),
	.A(\ab[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_4 (
	.S(\SUMB[7][4] ),
	.CO(\CARRYB[7][4] ),
	.CI(\SUMB[6][5] ),
	.B(\CARRYB[6][4] ),
	.A(\ab[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_3 (
	.S(\SUMB[7][3] ),
	.CO(\CARRYB[7][3] ),
	.CI(\SUMB[6][4] ),
	.B(\CARRYB[6][3] ),
	.A(\ab[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_2 (
	.S(\SUMB[7][2] ),
	.CO(\CARRYB[7][2] ),
	.CI(\SUMB[6][3] ),
	.B(\CARRYB[6][2] ),
	.A(\ab[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_1 (
	.S(\SUMB[7][1] ),
	.CO(\CARRYB[7][1] ),
	.CI(\SUMB[6][2] ),
	.B(\CARRYB[6][1] ),
	.A(\ab[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U2 (
	.Y(n3),
	.B(\ab[1][5] ),
	.A(\ab[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U3 (
	.Y(n4),
	.B(\ab[1][4] ),
	.A(\ab[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U4 (
	.Y(n5),
	.B(\ab[1][3] ),
	.A(\ab[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U5 (
	.Y(n6),
	.B(\ab[1][2] ),
	.A(\ab[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U6 (
	.Y(n7),
	.B(\ab[1][1] ),
	.A(\ab[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U7 (
	.Y(n8),
	.B(\ab[1][6] ),
	.A(\ab[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U8 (
	.Y(n9),
	.B(\ab[1][0] ),
	.A(\ab[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U9 (
	.Y(n10),
	.B(\ab[7][7] ),
	.A(\CARRYB[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U10 (
	.Y(n22),
	.A(\ab[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U11 (
	.Y(\A1[7] ),
	.B(\SUMB[7][2] ),
	.A(\CARRYB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U12 (
	.Y(PRODUCT[1]),
	.B(\ab[0][1] ),
	.A(\ab[1][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U13 (
	.Y(\A1[12] ),
	.B(\ab[7][7] ),
	.A(\CARRYB[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U14 (
	.Y(\A1[8] ),
	.B(\SUMB[7][3] ),
	.A(\CARRYB[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U15 (
	.Y(\A1[10] ),
	.B(\SUMB[7][5] ),
	.A(\CARRYB[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U16 (
	.Y(\A1[9] ),
	.B(\SUMB[7][4] ),
	.A(\CARRYB[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U17 (
	.Y(\A1[11] ),
	.B(\SUMB[7][6] ),
	.A(\CARRYB[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(n23),
	.A(\ab[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U19 (
	.Y(n21),
	.A(\ab[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n20),
	.A(\ab[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n19),
	.A(\ab[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n18),
	.A(\ab[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U23 (
	.Y(n11),
	.B(\SUMB[7][1] ),
	.A(\CARRYB[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U24 (
	.Y(n17),
	.A(\SUMB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U25 (
	.Y(n12),
	.B(\SUMB[7][2] ),
	.A(\CARRYB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U26 (
	.Y(n13),
	.B(\SUMB[7][4] ),
	.A(\CARRYB[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U27 (
	.Y(n14),
	.B(\SUMB[7][6] ),
	.A(\CARRYB[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U28 (
	.Y(n15),
	.B(\SUMB[7][3] ),
	.A(\CARRYB[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U29 (
	.Y(n16),
	.B(\SUMB[7][5] ),
	.A(\CARRYB[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U30 (
	.Y(\A1[6] ),
	.B(n17),
	.A(\CARRYB[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U31 (
	.Y(\SUMB[1][6] ),
	.B(n23),
	.A(\ab[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U32 (
	.Y(\SUMB[1][5] ),
	.B(n22),
	.A(\ab[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U33 (
	.Y(\SUMB[1][4] ),
	.B(n21),
	.A(\ab[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U34 (
	.Y(\SUMB[1][3] ),
	.B(n20),
	.A(\ab[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U35 (
	.Y(\SUMB[1][2] ),
	.B(n19),
	.A(\ab[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U36 (
	.Y(\SUMB[1][1] ),
	.B(n18),
	.A(\ab[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U37 (
	.Y(n32),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U38 (
	.Y(n33),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U39 (
	.Y(n38),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U40 (
	.Y(n39),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U41 (
	.Y(n36),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U42 (
	.Y(n37),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U43 (
	.Y(n34),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U44 (
	.Y(n35),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U45 (
	.Y(n25),
	.A(B[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U46 (
	.Y(n31),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U47 (
	.Y(n29),
	.A(B[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U48 (
	.Y(n28),
	.A(B[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U49 (
	.Y(n24),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U50 (
	.Y(n27),
	.A(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U51 (
	.Y(n26),
	.A(B[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U52 (
	.Y(n30),
	.A(B[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U54 (
	.Y(\ab[7][7] ),
	.B(n24),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U55 (
	.Y(\ab[7][6] ),
	.B(n25),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U56 (
	.Y(\ab[7][5] ),
	.B(n26),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U57 (
	.Y(\ab[7][4] ),
	.B(n27),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U58 (
	.Y(\ab[7][3] ),
	.B(n28),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U59 (
	.Y(\ab[7][2] ),
	.B(n29),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U60 (
	.Y(\ab[7][1] ),
	.B(n30),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U61 (
	.Y(\ab[7][0] ),
	.B(n31),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U62 (
	.Y(\ab[6][7] ),
	.B(n33),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U63 (
	.Y(\ab[6][6] ),
	.B(n33),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U64 (
	.Y(\ab[6][5] ),
	.B(n33),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U65 (
	.Y(\ab[6][4] ),
	.B(n33),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U66 (
	.Y(\ab[6][3] ),
	.B(n33),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U67 (
	.Y(\ab[6][2] ),
	.B(n33),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U68 (
	.Y(\ab[6][1] ),
	.B(n33),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U69 (
	.Y(\ab[6][0] ),
	.B(n33),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U70 (
	.Y(\ab[5][7] ),
	.B(n34),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U71 (
	.Y(\ab[5][6] ),
	.B(n34),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U72 (
	.Y(\ab[5][5] ),
	.B(n34),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U73 (
	.Y(\ab[5][4] ),
	.B(n34),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U74 (
	.Y(\ab[5][3] ),
	.B(n34),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U75 (
	.Y(\ab[5][2] ),
	.B(n34),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U76 (
	.Y(\ab[5][1] ),
	.B(n34),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U77 (
	.Y(\ab[5][0] ),
	.B(n34),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U78 (
	.Y(\ab[4][7] ),
	.B(n35),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U79 (
	.Y(\ab[4][6] ),
	.B(n35),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U80 (
	.Y(\ab[4][5] ),
	.B(n35),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U81 (
	.Y(\ab[4][4] ),
	.B(n35),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U82 (
	.Y(\ab[4][3] ),
	.B(n35),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U83 (
	.Y(\ab[4][2] ),
	.B(n35),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U84 (
	.Y(\ab[4][1] ),
	.B(n35),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U85 (
	.Y(\ab[4][0] ),
	.B(n35),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U86 (
	.Y(\ab[3][7] ),
	.B(n36),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U87 (
	.Y(\ab[3][6] ),
	.B(n36),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U88 (
	.Y(\ab[3][5] ),
	.B(n36),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U89 (
	.Y(\ab[3][4] ),
	.B(n36),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U90 (
	.Y(\ab[3][3] ),
	.B(n36),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U91 (
	.Y(\ab[3][2] ),
	.B(n36),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U92 (
	.Y(\ab[3][1] ),
	.B(n36),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U93 (
	.Y(\ab[3][0] ),
	.B(n36),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U94 (
	.Y(\ab[2][7] ),
	.B(n37),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U95 (
	.Y(\ab[2][6] ),
	.B(n37),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U96 (
	.Y(\ab[2][5] ),
	.B(n37),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U97 (
	.Y(\ab[2][4] ),
	.B(n37),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U98 (
	.Y(\ab[2][3] ),
	.B(n37),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U99 (
	.Y(\ab[2][2] ),
	.B(n37),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U100 (
	.Y(\ab[2][1] ),
	.B(n37),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U101 (
	.Y(\ab[2][0] ),
	.B(n37),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U102 (
	.Y(\ab[1][7] ),
	.B(n38),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U103 (
	.Y(\ab[1][6] ),
	.B(n38),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U104 (
	.Y(\ab[1][5] ),
	.B(n38),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U105 (
	.Y(\ab[1][4] ),
	.B(n38),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U106 (
	.Y(\ab[1][3] ),
	.B(n38),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U107 (
	.Y(\ab[1][2] ),
	.B(n38),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U108 (
	.Y(\ab[1][1] ),
	.B(n38),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U109 (
	.Y(\ab[1][0] ),
	.B(n38),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U110 (
	.Y(\ab[0][7] ),
	.B(n39),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U111 (
	.Y(\ab[0][6] ),
	.B(n39),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U112 (
	.Y(\ab[0][5] ),
	.B(n39),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U113 (
	.Y(\ab[0][4] ),
	.B(n39),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U114 (
	.Y(\ab[0][3] ),
	.B(n39),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U115 (
	.Y(\ab[0][2] ),
	.B(n39),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U116 (
	.Y(\ab[0][1] ),
	.B(n39),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U117 (
	.Y(PRODUCT[0]),
	.B(n39),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_RTL_DATA_WIDTH8_DW01_add_1 FS_1 (
	.A({ 1'b0,
		\A1[12] ,
		\A1[11] ,
		\A1[10] ,
		\A1[9] ,
		\A1[8] ,
		\A1[7] ,
		\A1[6] ,
		\SUMB[7][0] ,
		\A1[4] ,
		\A1[3] ,
		\A1[2] ,
		\A1[1] ,
		\A1[0]  }),
	.B({ n10,
		n14,
		n16,
		n13,
		n15,
		n12,
		n11,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0 }),
	.CI(1'b0),
	.SUM({ PRODUCT[15],
		PRODUCT[14],
		PRODUCT[13],
		PRODUCT[12],
		PRODUCT[11],
		PRODUCT[10],
		PRODUCT[9],
		PRODUCT[8],
		PRODUCT[7],
		PRODUCT[6],
		PRODUCT[5],
		PRODUCT[4],
		PRODUCT[3],
		PRODUCT[2] }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_RTL_DATA_WIDTH8_DW01_add_1 (
	A, 
	B, 
	CI, 
	SUM, 
	CO, 
	VDD, 
	VSS);
   input [13:0] A;
   input [13:0] B;
   input CI;
   output [13:0] SUM;
   output CO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \A[5] ;
   wire \A[4] ;
   wire \A[3] ;
   wire \A[2] ;
   wire \A[1] ;
   wire \A[0] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;

   assign SUM[6] = A[6] ;
   assign SUM[5] = \A[5]  ;
   assign \A[5]  = A[5] ;
   assign SUM[4] = \A[4]  ;
   assign \A[4]  = A[4] ;
   assign SUM[3] = \A[3]  ;
   assign \A[3]  = A[3] ;
   assign SUM[2] = \A[2]  ;
   assign \A[2]  = A[2] ;
   assign SUM[1] = \A[1]  ;
   assign \A[1]  = A[1] ;
   assign SUM[0] = \A[0]  ;
   assign \A[0]  = A[0] ;

   // Module instantiations
   AOI21BX2M U2 (
	.Y(n1),
	.B0N(n12),
	.A1(A[12]),
	.A0(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U3 (
	.Y(n8),
	.B(B[7]),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U4 (
	.Y(SUM[7]),
	.B(n2),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(n2),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U6 (
	.Y(SUM[13]),
	.B(n1),
	.A(B[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U7 (
	.Y(SUM[9]),
	.B(n4),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U8 (
	.Y(n4),
	.B(n6),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U9 (
	.Y(SUM[8]),
	.B(n8),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U10 (
	.Y(n7),
	.B(n10),
	.AN(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U11 (
	.Y(n12),
	.B0(B[12]),
	.A1(n11),
	.A0(A[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U12 (
	.Y(SUM[12]),
	.C(n11),
	.B(A[12]),
	.A(B[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21BX1M U13 (
	.Y(n11),
	.B0N(n15),
	.A1(n14),
	.A0(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U14 (
	.Y(SUM[11]),
	.B(n16),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U15 (
	.Y(n16),
	.B(n13),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U16 (
	.Y(n13),
	.B(A[11]),
	.A(B[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U17 (
	.Y(n15),
	.B(A[11]),
	.A(B[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U18 (
	.Y(n14),
	.B0(n19),
	.A1(n18),
	.A0(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U19 (
	.Y(SUM[10]),
	.B(n18),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X1M U20 (
	.Y(n18),
	.B0(n5),
	.A1N(n6),
	.A0N(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U21 (
	.Y(n5),
	.B(A[9]),
	.A(B[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U22 (
	.Y(n6),
	.B(A[9]),
	.A(B[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U23 (
	.Y(n3),
	.B0(n10),
	.A1(n9),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U24 (
	.Y(n10),
	.B(A[8]),
	.A(B[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U25 (
	.Y(n9),
	.B(A[8]),
	.A(B[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U26 (
	.Y(n20),
	.B(n19),
	.AN(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U27 (
	.Y(n19),
	.B(A[10]),
	.A(B[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U28 (
	.Y(n17),
	.B(A[10]),
	.A(B[10]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_TOP_DATA_WIDTH_TOP8_FIFO_DEPTH_TOP8_ADDRESS_BITS_TOP3_test_1 (
	W_CLK, 
	W_RST, 
	R_CLK, 
	R_RST, 
	WINC, 
	RINC, 
	W_DATA, 
	W_FULL, 
	R_EMPTY, 
	R_DATA, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN13_SE, 
	FE_OFN5_scanclkref__L2_N0, 
	VDD, 
	VSS);
   input W_CLK;
   input W_RST;
   input R_CLK;
   input R_RST;
   input WINC;
   input RINC;
   input [7:0] W_DATA;
   output W_FULL;
   output R_EMPTY;
   output [7:0] R_DATA;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN13_SE;
   input FE_OFN5_scanclkref__L2_N0;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN6_scanclkref__L1_N0;
   wire FE_OFN15_SE;
   wire FE_OFN6_scanclkref;
   wire FE_OFN2_scanrst2;
   wire n5;
   wire [2:0] W_ADDRESS;
   wire [2:0] R_ADDRESS;
   wire [3:0] WQ2_RPTR;
   wire [3:0] W_PTR;
   wire [3:0] RQ2_WPTR;
   wire [3:0] R_PTR;

   assign test_so = W_PTR[3] ;

   // Module instantiations
   CLKBUFX40M FE_OFN6_scanclkref__L1_I0 (
	.Y(FE_OFN6_scanclkref__L1_N0),
	.A(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX4M FE_OFC15_SE (
	.Y(FE_OFN15_SE),
	.A(FE_OFN13_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX8M FE_OFC6_scanclkref (
	.Y(FE_OFN6_scanclkref),
	.A(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX8M FE_OFC2_scanrst2 (
	.Y(FE_OFN2_scanrst2),
	.A(W_RST), 
	.VDD(VDD), 
	.VSS(VSS));
   FIFO_BUFFER_DATA_WIDTH8_FIFO_DEPTH8_ADDRESS_BITS3_test_1 FIFO_BUFFER (
	.W_CLK(FE_OFN5_scanclkref__L2_N0),
	.W_RST(W_RST),
	.WINC(WINC),
	.W_FULL(W_FULL),
	.W_DATA({ W_DATA[7],
		W_DATA[6],
		W_DATA[5],
		W_DATA[4],
		W_DATA[3],
		W_DATA[2],
		W_DATA[1],
		W_DATA[0] }),
	.W_ADDRESS({ W_ADDRESS[2],
		W_ADDRESS[1],
		W_ADDRESS[0] }),
	.R_ADDRESS({ R_ADDRESS[2],
		R_ADDRESS[1],
		R_ADDRESS[0] }),
	.R_DATA({ R_DATA[7],
		R_DATA[6],
		R_DATA[5],
		R_DATA[4],
		R_DATA[3],
		R_DATA[2],
		R_DATA[1],
		R_DATA[0] }),
	.test_si(n5),
	.test_se(test_se),
	.FE_OFN2_scanrst2(FE_OFN2_scanrst2),
	.FE_OFN6_scanclkref(FE_OFN6_scanclkref__L1_N0),
	.FE_OFN13_SE(FE_OFN13_SE),
	.FE_OFN15_SE(FE_OFN15_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   FIFO_WR_ADDRESS_BITS3_test_1 FIFO_WR (
	.W_CLK(FE_OFN5_scanclkref__L2_N0),
	.W_RST(W_RST),
	.WINC(WINC),
	.RINC(RINC),
	.WQ2_RPTR({ WQ2_RPTR[3],
		WQ2_RPTR[2],
		WQ2_RPTR[1],
		WQ2_RPTR[0] }),
	.W_FULL(W_FULL),
	.W_ADDRESS({ W_ADDRESS[2],
		W_ADDRESS[1],
		W_ADDRESS[0] }),
	.W_PTR({ W_PTR[3],
		W_PTR[2],
		W_PTR[1],
		W_PTR[0] }),
	.test_si(R_PTR[3]),
	.test_se(test_se),
	.FE_OFN6_scanclkref(FE_OFN6_scanclkref__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   FIFO_RD_ADDRESS_BITS3_test_1 FIFO_RD (
	.R_CLK(R_CLK),
	.R_RST(R_RST),
	.RINC(RINC),
	.RQ2_WPTR({ RQ2_WPTR[3],
		RQ2_WPTR[2],
		RQ2_WPTR[1],
		RQ2_WPTR[0] }),
	.R_EMPTY(R_EMPTY),
	.R_ADDRESS({ R_ADDRESS[2],
		R_ADDRESS[1],
		R_ADDRESS[0] }),
	.R_PTR({ R_PTR[3],
		R_PTR[2],
		R_PTR[1],
		R_PTR[0] }),
	.test_si(R_DATA[7]),
	.test_se(FE_OFN13_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   DF_SYNC_ADDRESS_BITS3_test_1 DF_SYNC (
	.W_CLK(FE_OFN5_scanclkref__L2_N0),
	.W_RST(FE_OFN2_scanrst2),
	.R_CLK(R_CLK),
	.R_RST(R_RST),
	.W_PTR({ W_PTR[3],
		W_PTR[2],
		W_PTR[1],
		W_PTR[0] }),
	.R_PTR({ R_PTR[3],
		R_PTR[2],
		R_PTR[1],
		R_PTR[0] }),
	.RQ2_WPTR({ RQ2_WPTR[3],
		RQ2_WPTR[2],
		RQ2_WPTR[1],
		RQ2_WPTR[0] }),
	.WQ2_RPTR({ WQ2_RPTR[3],
		WQ2_RPTR[2],
		WQ2_RPTR[1],
		WQ2_RPTR[0] }),
	.test_si(test_si),
	.test_so(n5),
	.test_se(FE_OFN13_SE),
	.FE_OFN15_SE(FE_OFN15_SE), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_BUFFER_DATA_WIDTH8_FIFO_DEPTH8_ADDRESS_BITS3_test_1 (
	W_CLK, 
	W_RST, 
	WINC, 
	W_FULL, 
	W_DATA, 
	W_ADDRESS, 
	R_ADDRESS, 
	R_DATA, 
	test_si, 
	test_se, 
	FE_OFN2_scanrst2, 
	FE_OFN6_scanclkref, 
	FE_OFN13_SE, 
	FE_OFN15_SE, 
	VDD, 
	VSS);
   input W_CLK;
   input W_RST;
   input WINC;
   input W_FULL;
   input [7:0] W_DATA;
   input [2:0] W_ADDRESS;
   input [2:0] R_ADDRESS;
   output [7:0] R_DATA;
   input test_si;
   input test_se;
   input FE_OFN2_scanrst2;
   input FE_OFN6_scanclkref;
   input FE_OFN13_SE;
   input FE_OFN15_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N9;
   wire N10;
   wire N11;
   wire \REG[7][7] ;
   wire \REG[7][6] ;
   wire \REG[7][5] ;
   wire \REG[7][4] ;
   wire \REG[7][3] ;
   wire \REG[7][2] ;
   wire \REG[7][1] ;
   wire \REG[7][0] ;
   wire \REG[6][7] ;
   wire \REG[6][6] ;
   wire \REG[6][5] ;
   wire \REG[6][4] ;
   wire \REG[6][3] ;
   wire \REG[6][2] ;
   wire \REG[6][1] ;
   wire \REG[6][0] ;
   wire \REG[5][7] ;
   wire \REG[5][6] ;
   wire \REG[5][5] ;
   wire \REG[5][4] ;
   wire \REG[5][3] ;
   wire \REG[5][2] ;
   wire \REG[5][1] ;
   wire \REG[5][0] ;
   wire \REG[4][7] ;
   wire \REG[4][6] ;
   wire \REG[4][5] ;
   wire \REG[4][4] ;
   wire \REG[4][3] ;
   wire \REG[4][2] ;
   wire \REG[4][1] ;
   wire \REG[4][0] ;
   wire \REG[3][7] ;
   wire \REG[3][6] ;
   wire \REG[3][5] ;
   wire \REG[3][4] ;
   wire \REG[3][3] ;
   wire \REG[3][2] ;
   wire \REG[3][1] ;
   wire \REG[3][0] ;
   wire \REG[2][7] ;
   wire \REG[2][6] ;
   wire \REG[2][5] ;
   wire \REG[2][4] ;
   wire \REG[2][3] ;
   wire \REG[2][2] ;
   wire \REG[2][1] ;
   wire \REG[2][0] ;
   wire \REG[1][7] ;
   wire \REG[1][6] ;
   wire \REG[1][5] ;
   wire \REG[1][4] ;
   wire \REG[1][3] ;
   wire \REG[1][2] ;
   wire \REG[1][1] ;
   wire \REG[1][0] ;
   wire \REG[0][7] ;
   wire \REG[0][6] ;
   wire \REG[0][5] ;
   wire \REG[0][4] ;
   wire \REG[0][3] ;
   wire \REG[0][2] ;
   wire \REG[0][1] ;
   wire \REG[0][0] ;
   wire N31;
   wire N32;
   wire N33;
   wire N34;
   wire N35;
   wire N36;
   wire N37;
   wire N38;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;

   assign N9 = R_ADDRESS[0] ;
   assign N10 = R_ADDRESS[1] ;
   assign N11 = R_ADDRESS[2] ;

   // Module instantiations
   SDFFRQX2M \REG_reg[5][7]  (
	.SI(\REG[5][6] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[5][7] ),
	.D(n141),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[5][6]  (
	.SI(\REG[5][5] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[5][6] ),
	.D(n140),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[5][5]  (
	.SI(\REG[5][4] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[5][5] ),
	.D(n139),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[5][4]  (
	.SI(\REG[5][3] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[5][4] ),
	.D(n138),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[5][3]  (
	.SI(\REG[5][2] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[5][3] ),
	.D(n137),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[5][2]  (
	.SI(\REG[5][1] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[5][2] ),
	.D(n136),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[5][1]  (
	.SI(\REG[5][0] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[5][1] ),
	.D(n135),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[5][0]  (
	.SI(\REG[4][7] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[5][0] ),
	.D(n134),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[1][7]  (
	.SI(\REG[1][6] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[1][7] ),
	.D(n109),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[1][6]  (
	.SI(\REG[1][5] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[1][6] ),
	.D(n108),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[1][5]  (
	.SI(\REG[1][4] ),
	.SE(FE_OFN15_SE),
	.RN(W_RST),
	.Q(\REG[1][5] ),
	.D(n107),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[1][4]  (
	.SI(\REG[1][3] ),
	.SE(test_se),
	.RN(W_RST),
	.Q(\REG[1][4] ),
	.D(n106),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[1][3]  (
	.SI(\REG[1][2] ),
	.SE(FE_OFN15_SE),
	.RN(W_RST),
	.Q(\REG[1][3] ),
	.D(n105),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[1][2]  (
	.SI(\REG[1][1] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[1][2] ),
	.D(n104),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[1][1]  (
	.SI(\REG[1][0] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[1][1] ),
	.D(n103),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[1][0]  (
	.SI(\REG[0][7] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[1][0] ),
	.D(n102),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[7][7]  (
	.SI(\REG[7][6] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[7][7] ),
	.D(n157),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[7][6]  (
	.SI(\REG[7][5] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[7][6] ),
	.D(n156),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[7][5]  (
	.SI(\REG[7][4] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[7][5] ),
	.D(n155),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[7][4]  (
	.SI(\REG[7][3] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[7][4] ),
	.D(n154),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[7][3]  (
	.SI(\REG[7][2] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[7][3] ),
	.D(n153),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[7][2]  (
	.SI(\REG[7][1] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[7][2] ),
	.D(n152),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[7][1]  (
	.SI(\REG[7][0] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[7][1] ),
	.D(n151),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[7][0]  (
	.SI(\REG[6][7] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[7][0] ),
	.D(n150),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[3][7]  (
	.SI(\REG[3][6] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[3][7] ),
	.D(n125),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[3][6]  (
	.SI(\REG[3][5] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[3][6] ),
	.D(n124),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[3][5]  (
	.SI(\REG[3][4] ),
	.SE(FE_OFN15_SE),
	.RN(W_RST),
	.Q(\REG[3][5] ),
	.D(n123),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[3][4]  (
	.SI(\REG[3][3] ),
	.SE(FE_OFN15_SE),
	.RN(W_RST),
	.Q(\REG[3][4] ),
	.D(n122),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[3][3]  (
	.SI(\REG[3][2] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[3][3] ),
	.D(n121),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[3][2]  (
	.SI(\REG[3][1] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[3][2] ),
	.D(n120),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[3][1]  (
	.SI(\REG[3][0] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[3][1] ),
	.D(n119),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[3][0]  (
	.SI(\REG[2][7] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[3][0] ),
	.D(n118),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[6][7]  (
	.SI(\REG[6][6] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[6][7] ),
	.D(n149),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[6][6]  (
	.SI(\REG[6][5] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[6][6] ),
	.D(n148),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[6][5]  (
	.SI(\REG[6][4] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[6][5] ),
	.D(n147),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[6][4]  (
	.SI(\REG[6][3] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[6][4] ),
	.D(n146),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[6][3]  (
	.SI(\REG[6][2] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[6][3] ),
	.D(n145),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[6][2]  (
	.SI(\REG[6][1] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[6][2] ),
	.D(n144),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[6][1]  (
	.SI(\REG[6][0] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[6][1] ),
	.D(n143),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[6][0]  (
	.SI(\REG[5][7] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[6][0] ),
	.D(n142),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[2][7]  (
	.SI(\REG[2][6] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[2][7] ),
	.D(n117),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[2][6]  (
	.SI(\REG[2][5] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[2][6] ),
	.D(n116),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[2][5]  (
	.SI(\REG[2][4] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[2][5] ),
	.D(n115),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[2][4]  (
	.SI(\REG[2][3] ),
	.SE(FE_OFN15_SE),
	.RN(W_RST),
	.Q(\REG[2][4] ),
	.D(n114),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[2][3]  (
	.SI(\REG[2][2] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[2][3] ),
	.D(n113),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[2][2]  (
	.SI(\REG[2][1] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[2][2] ),
	.D(n112),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[2][1]  (
	.SI(\REG[2][0] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[2][1] ),
	.D(n111),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[2][0]  (
	.SI(\REG[1][7] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[2][0] ),
	.D(n110),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[4][7]  (
	.SI(\REG[4][6] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[4][7] ),
	.D(n133),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[4][6]  (
	.SI(\REG[4][5] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[4][6] ),
	.D(n132),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[4][5]  (
	.SI(\REG[4][4] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[4][5] ),
	.D(n131),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[4][4]  (
	.SI(\REG[4][3] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[4][4] ),
	.D(n130),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[4][3]  (
	.SI(\REG[4][2] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[4][3] ),
	.D(n129),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[4][2]  (
	.SI(\REG[4][1] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[4][2] ),
	.D(n128),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[4][1]  (
	.SI(\REG[4][0] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[4][1] ),
	.D(n127),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[4][0]  (
	.SI(\REG[3][7] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[4][0] ),
	.D(n126),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0][7]  (
	.SI(\REG[0][6] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[0][7] ),
	.D(n101),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0][6]  (
	.SI(\REG[0][5] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[0][6] ),
	.D(n100),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0][5]  (
	.SI(\REG[0][4] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[0][5] ),
	.D(n99),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0][4]  (
	.SI(\REG[0][3] ),
	.SE(test_se),
	.RN(W_RST),
	.Q(\REG[0][4] ),
	.D(n98),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0][3]  (
	.SI(\REG[0][2] ),
	.SE(FE_OFN15_SE),
	.RN(W_RST),
	.Q(\REG[0][3] ),
	.D(n97),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0][2]  (
	.SI(\REG[0][1] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[0][2] ),
	.D(n96),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0][1]  (
	.SI(\REG[0][0] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[0][1] ),
	.D(n95),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0][0]  (
	.SI(test_si),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(\REG[0][0] ),
	.D(n94),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R_DATA_reg[5]  (
	.SI(R_DATA[4]),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(R_DATA[5]),
	.D(N33),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R_DATA_reg[1]  (
	.SI(R_DATA[0]),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(R_DATA[1]),
	.D(N37),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R_DATA_reg[4]  (
	.SI(R_DATA[3]),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(R_DATA[4]),
	.D(N34),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R_DATA_reg[0]  (
	.SI(\REG[7][7] ),
	.SE(FE_OFN15_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(R_DATA[0]),
	.D(N38),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R_DATA_reg[3]  (
	.SI(R_DATA[2]),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(R_DATA[3]),
	.D(N35),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R_DATA_reg[2]  (
	.SI(R_DATA[1]),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(R_DATA[2]),
	.D(N36),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R_DATA_reg[6]  (
	.SI(R_DATA[5]),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(R_DATA[6]),
	.D(N32),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R_DATA_reg[7]  (
	.SI(R_DATA[6]),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_scanrst2),
	.Q(R_DATA[7]),
	.D(N31),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U92 (
	.Y(n91),
	.B(W_FULL),
	.AN(WINC), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U97 (
	.Y(n92),
	.C(n85),
	.B(n187),
	.A(n186), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U98 (
	.Y(n86),
	.C(n87),
	.B(n187),
	.A(n186), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U99 (
	.Y(n93),
	.C(W_ADDRESS[0]),
	.B(n187),
	.A(n85), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U100 (
	.Y(n85),
	.B(W_ADDRESS[2]),
	.AN(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U101 (
	.Y(n187),
	.A(W_ADDRESS[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U102 (
	.Y(n186),
	.A(W_ADDRESS[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U103 (
	.Y(n102),
	.B1(n93),
	.B0(n195),
	.A1N(n93),
	.A0N(\REG[1][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U104 (
	.Y(n103),
	.B1(n93),
	.B0(n194),
	.A1N(n93),
	.A0N(\REG[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U105 (
	.Y(n104),
	.B1(n93),
	.B0(n193),
	.A1N(n93),
	.A0N(\REG[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U106 (
	.Y(n105),
	.B1(n93),
	.B0(n192),
	.A1N(n93),
	.A0N(\REG[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U107 (
	.Y(n106),
	.B1(n93),
	.B0(n191),
	.A1N(n93),
	.A0N(\REG[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U108 (
	.Y(n107),
	.B1(n93),
	.B0(n190),
	.A1N(n93),
	.A0N(\REG[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U109 (
	.Y(n108),
	.B1(n93),
	.B0(n189),
	.A1N(n93),
	.A0N(\REG[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U110 (
	.Y(n109),
	.B1(n93),
	.B0(n188),
	.A1N(n93),
	.A0N(\REG[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U111 (
	.Y(n94),
	.B1(n92),
	.B0(n195),
	.A1N(n92),
	.A0N(\REG[0][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U112 (
	.Y(n95),
	.B1(n92),
	.B0(n194),
	.A1N(n92),
	.A0N(\REG[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U113 (
	.Y(n96),
	.B1(n92),
	.B0(n193),
	.A1N(n92),
	.A0N(\REG[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U114 (
	.Y(n97),
	.B1(n92),
	.B0(n192),
	.A1N(n92),
	.A0N(\REG[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U115 (
	.Y(n98),
	.B1(n92),
	.B0(n191),
	.A1N(n92),
	.A0N(\REG[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U116 (
	.Y(n99),
	.B1(n92),
	.B0(n190),
	.A1N(n92),
	.A0N(\REG[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U117 (
	.Y(n100),
	.B1(n92),
	.B0(n189),
	.A1N(n92),
	.A0N(\REG[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U118 (
	.Y(n101),
	.B1(n92),
	.B0(n188),
	.A1N(n92),
	.A0N(\REG[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U119 (
	.Y(n126),
	.B1(n86),
	.B0(n195),
	.A1N(n86),
	.A0N(\REG[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U120 (
	.Y(n127),
	.B1(n86),
	.B0(n194),
	.A1N(n86),
	.A0N(\REG[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U121 (
	.Y(n128),
	.B1(n86),
	.B0(n193),
	.A1N(n86),
	.A0N(\REG[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U122 (
	.Y(n129),
	.B1(n86),
	.B0(n192),
	.A1N(n86),
	.A0N(\REG[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U123 (
	.Y(n130),
	.B1(n86),
	.B0(n191),
	.A1N(n86),
	.A0N(\REG[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U124 (
	.Y(n131),
	.B1(n86),
	.B0(n190),
	.A1N(n86),
	.A0N(\REG[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U125 (
	.Y(n132),
	.B1(n86),
	.B0(n189),
	.A1N(n86),
	.A0N(\REG[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U126 (
	.Y(n133),
	.B1(n86),
	.B0(n188),
	.A1N(n86),
	.A0N(\REG[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX4M U127 (
	.Y(n164),
	.A(N9), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U128 (
	.Y(n195),
	.A(W_DATA[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U129 (
	.Y(n194),
	.A(W_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U130 (
	.Y(n193),
	.A(W_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U131 (
	.Y(n192),
	.A(W_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U132 (
	.Y(n191),
	.A(W_DATA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U133 (
	.Y(n190),
	.A(W_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U134 (
	.Y(n189),
	.A(W_DATA[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U135 (
	.Y(n188),
	.A(W_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U136 (
	.Y(n123),
	.B1(n84),
	.B0(n190),
	.A1N(n84),
	.A0N(\REG[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U137 (
	.Y(n124),
	.B1(n84),
	.B0(n189),
	.A1N(n84),
	.A0N(\REG[3][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U138 (
	.Y(n125),
	.B1(n84),
	.B0(n188),
	.A1N(n84),
	.A0N(\REG[3][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U139 (
	.Y(n134),
	.B1(n88),
	.B0(n195),
	.A1N(n88),
	.A0N(\REG[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U140 (
	.Y(n135),
	.B1(n88),
	.B0(n194),
	.A1N(n88),
	.A0N(\REG[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U141 (
	.Y(n136),
	.B1(n88),
	.B0(n193),
	.A1N(n88),
	.A0N(\REG[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U142 (
	.Y(n137),
	.B1(n88),
	.B0(n192),
	.A1N(n88),
	.A0N(\REG[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U143 (
	.Y(n138),
	.B1(n88),
	.B0(n191),
	.A1N(n88),
	.A0N(\REG[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U144 (
	.Y(n139),
	.B1(n88),
	.B0(n190),
	.A1N(n88),
	.A0N(\REG[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U145 (
	.Y(n140),
	.B1(n88),
	.B0(n189),
	.A1N(n88),
	.A0N(\REG[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U146 (
	.Y(n141),
	.B1(n88),
	.B0(n188),
	.A1N(n88),
	.A0N(\REG[5][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U147 (
	.Y(n142),
	.B1(n89),
	.B0(n195),
	.A1N(n89),
	.A0N(\REG[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U148 (
	.Y(n143),
	.B1(n89),
	.B0(n194),
	.A1N(n89),
	.A0N(\REG[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U149 (
	.Y(n144),
	.B1(n89),
	.B0(n193),
	.A1N(n89),
	.A0N(\REG[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U150 (
	.Y(n145),
	.B1(n89),
	.B0(n192),
	.A1N(n89),
	.A0N(\REG[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U151 (
	.Y(n146),
	.B1(n89),
	.B0(n191),
	.A1N(n89),
	.A0N(\REG[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U152 (
	.Y(n147),
	.B1(n89),
	.B0(n190),
	.A1N(n89),
	.A0N(\REG[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U153 (
	.Y(n148),
	.B1(n89),
	.B0(n189),
	.A1N(n89),
	.A0N(\REG[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U154 (
	.Y(n149),
	.B1(n89),
	.B0(n188),
	.A1N(n89),
	.A0N(\REG[6][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U155 (
	.Y(n150),
	.B1(n90),
	.B0(n195),
	.A1N(n90),
	.A0N(\REG[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U156 (
	.Y(n151),
	.B1(n90),
	.B0(n194),
	.A1N(n90),
	.A0N(\REG[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U157 (
	.Y(n152),
	.B1(n90),
	.B0(n193),
	.A1N(n90),
	.A0N(\REG[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U158 (
	.Y(n153),
	.B1(n90),
	.B0(n192),
	.A1N(n90),
	.A0N(\REG[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U159 (
	.Y(n154),
	.B1(n90),
	.B0(n191),
	.A1N(n90),
	.A0N(\REG[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U160 (
	.Y(n155),
	.B1(n90),
	.B0(n190),
	.A1N(n90),
	.A0N(\REG[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U161 (
	.Y(n156),
	.B1(n90),
	.B0(n189),
	.A1N(n90),
	.A0N(\REG[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U162 (
	.Y(n157),
	.B1(n90),
	.B0(n188),
	.A1N(n90),
	.A0N(\REG[7][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U163 (
	.Y(n110),
	.B1(n195),
	.B0(n83),
	.A1N(n83),
	.A0N(\REG[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U164 (
	.Y(n111),
	.B1(n194),
	.B0(n83),
	.A1N(n83),
	.A0N(\REG[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U165 (
	.Y(n112),
	.B1(n193),
	.B0(n83),
	.A1N(n83),
	.A0N(\REG[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U166 (
	.Y(n113),
	.B1(n192),
	.B0(n83),
	.A1N(n83),
	.A0N(\REG[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U167 (
	.Y(n114),
	.B1(n191),
	.B0(n83),
	.A1N(n83),
	.A0N(\REG[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U168 (
	.Y(n115),
	.B1(n190),
	.B0(n83),
	.A1N(n83),
	.A0N(\REG[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U169 (
	.Y(n116),
	.B1(n189),
	.B0(n83),
	.A1N(n83),
	.A0N(\REG[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U170 (
	.Y(n117),
	.B1(n188),
	.B0(n83),
	.A1N(n83),
	.A0N(\REG[2][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U171 (
	.Y(n118),
	.B1(n195),
	.B0(n84),
	.A1N(n84),
	.A0N(\REG[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U172 (
	.Y(n119),
	.B1(n194),
	.B0(n84),
	.A1N(n84),
	.A0N(\REG[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U173 (
	.Y(n120),
	.B1(n193),
	.B0(n84),
	.A1N(n84),
	.A0N(\REG[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U174 (
	.Y(n121),
	.B1(n192),
	.B0(n84),
	.A1N(n84),
	.A0N(\REG[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U175 (
	.Y(n122),
	.B1(n191),
	.B0(n84),
	.A1N(n84),
	.A0N(\REG[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U176 (
	.Y(n87),
	.B(n91),
	.A(W_ADDRESS[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U177 (
	.Y(n90),
	.C(n87),
	.B(W_ADDRESS[1]),
	.A(W_ADDRESS[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U178 (
	.Y(n89),
	.C(n87),
	.B(n186),
	.A(W_ADDRESS[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U179 (
	.Y(n88),
	.C(n87),
	.B(n187),
	.A(W_ADDRESS[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U180 (
	.Y(n84),
	.C(W_ADDRESS[0]),
	.B(n85),
	.A(W_ADDRESS[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U181 (
	.Y(n83),
	.C(W_ADDRESS[1]),
	.B(n186),
	.A(n85), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U182 (
	.Y(N38),
	.S0(N11),
	.B(n73),
	.A(n74), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U183 (
	.Y(n73),
	.S1(N10),
	.S0(n164),
	.D(\REG[7][0] ),
	.C(\REG[6][0] ),
	.B(\REG[5][0] ),
	.A(\REG[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U184 (
	.Y(n74),
	.S1(N10),
	.S0(n164),
	.D(\REG[3][0] ),
	.C(\REG[2][0] ),
	.B(\REG[1][0] ),
	.A(\REG[0][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U185 (
	.Y(N37),
	.S0(N11),
	.B(n75),
	.A(n76), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U186 (
	.Y(n75),
	.S1(N10),
	.S0(n164),
	.D(\REG[7][1] ),
	.C(\REG[6][1] ),
	.B(\REG[5][1] ),
	.A(\REG[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U187 (
	.Y(n76),
	.S1(N10),
	.S0(n164),
	.D(\REG[3][1] ),
	.C(\REG[2][1] ),
	.B(\REG[1][1] ),
	.A(\REG[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U188 (
	.Y(N36),
	.S0(N11),
	.B(n77),
	.A(n78), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U189 (
	.Y(n77),
	.S1(N10),
	.S0(n164),
	.D(\REG[7][2] ),
	.C(\REG[6][2] ),
	.B(\REG[5][2] ),
	.A(\REG[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U190 (
	.Y(n78),
	.S1(N10),
	.S0(n164),
	.D(\REG[3][2] ),
	.C(\REG[2][2] ),
	.B(\REG[1][2] ),
	.A(\REG[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U191 (
	.Y(N35),
	.S0(N11),
	.B(n79),
	.A(n80), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U192 (
	.Y(n79),
	.S1(N10),
	.S0(n164),
	.D(\REG[7][3] ),
	.C(\REG[6][3] ),
	.B(\REG[5][3] ),
	.A(\REG[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U193 (
	.Y(n80),
	.S1(N10),
	.S0(n164),
	.D(\REG[3][3] ),
	.C(\REG[2][3] ),
	.B(\REG[1][3] ),
	.A(\REG[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U194 (
	.Y(N34),
	.S0(N11),
	.B(n81),
	.A(n82), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U195 (
	.Y(n81),
	.S1(N10),
	.S0(n164),
	.D(\REG[7][4] ),
	.C(\REG[6][4] ),
	.B(\REG[5][4] ),
	.A(\REG[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U196 (
	.Y(n82),
	.S1(N10),
	.S0(n164),
	.D(\REG[3][4] ),
	.C(\REG[2][4] ),
	.B(\REG[1][4] ),
	.A(\REG[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U197 (
	.Y(N33),
	.S0(N11),
	.B(n158),
	.A(n159), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U198 (
	.Y(n158),
	.S1(N10),
	.S0(n164),
	.D(\REG[7][5] ),
	.C(\REG[6][5] ),
	.B(\REG[5][5] ),
	.A(\REG[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U199 (
	.Y(n159),
	.S1(N10),
	.S0(n164),
	.D(\REG[3][5] ),
	.C(\REG[2][5] ),
	.B(\REG[1][5] ),
	.A(\REG[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U200 (
	.Y(N32),
	.S0(N11),
	.B(n160),
	.A(n161), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U201 (
	.Y(n160),
	.S1(N10),
	.S0(n164),
	.D(\REG[7][6] ),
	.C(\REG[6][6] ),
	.B(\REG[5][6] ),
	.A(\REG[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U202 (
	.Y(n161),
	.S1(N10),
	.S0(n164),
	.D(\REG[3][6] ),
	.C(\REG[2][6] ),
	.B(\REG[1][6] ),
	.A(\REG[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U203 (
	.Y(N31),
	.S0(N11),
	.B(n162),
	.A(n163), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U204 (
	.Y(n162),
	.S1(N10),
	.S0(n164),
	.D(\REG[7][7] ),
	.C(\REG[6][7] ),
	.B(\REG[5][7] ),
	.A(\REG[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U205 (
	.Y(n163),
	.S1(N10),
	.S0(n164),
	.D(\REG[3][7] ),
	.C(\REG[2][7] ),
	.B(\REG[1][7] ),
	.A(\REG[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_WR_ADDRESS_BITS3_test_1 (
	W_CLK, 
	W_RST, 
	WINC, 
	RINC, 
	WQ2_RPTR, 
	W_FULL, 
	W_ADDRESS, 
	W_PTR, 
	test_si, 
	test_se, 
	FE_OFN6_scanclkref, 
	VDD, 
	VSS);
   input W_CLK;
   input W_RST;
   input WINC;
   input RINC;
   input [3:0] WQ2_RPTR;
   output W_FULL;
   output [2:0] W_ADDRESS;
   output [3:0] W_PTR;
   input test_si;
   input test_se;
   input FE_OFN6_scanclkref;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n12;
   wire n14;
   wire n16;
   wire n18;

   // Module instantiations
   SDFFRQX2M \add_ptr_reg[3]  (
	.SI(W_ADDRESS[2]),
	.SE(test_se),
	.RN(W_RST),
	.Q(W_PTR[3]),
	.D(n18),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \add_ptr_reg[2]  (
	.SI(W_ADDRESS[1]),
	.SE(test_se),
	.RN(W_RST),
	.Q(W_ADDRESS[2]),
	.D(n14),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \add_ptr_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(W_RST),
	.Q(W_ADDRESS[0]),
	.D(n16),
	.CK(FE_OFN6_scanclkref), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \add_ptr_reg[1]  (
	.SI(W_ADDRESS[0]),
	.SE(test_se),
	.RN(W_RST),
	.Q(W_ADDRESS[1]),
	.D(n12),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U3 (
	.Y(n3),
	.B(n4),
	.A(WINC), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U4 (
	.Y(W_FULL),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U5 (
	.Y(n1),
	.B(n3),
	.AN(W_ADDRESS[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U6 (
	.Y(n6),
	.B(WQ2_RPTR[0]),
	.A(W_PTR[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U7 (
	.Y(n18),
	.B(n5),
	.A(W_PTR[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U8 (
	.Y(n5),
	.C(n1),
	.B(W_ADDRESS[2]),
	.A(W_ADDRESS[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U9 (
	.Y(n16),
	.B(n3),
	.A(W_ADDRESS[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U10 (
	.Y(n14),
	.B(n2),
	.A(W_ADDRESS[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U11 (
	.Y(n2),
	.B(W_ADDRESS[1]),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U12 (
	.Y(n4),
	.D(n9),
	.C(n8),
	.B(n7),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U13 (
	.Y(n8),
	.B(W_PTR[2]),
	.A(WQ2_RPTR[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U14 (
	.Y(n9),
	.B(WQ2_RPTR[3]),
	.A(W_PTR[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U15 (
	.Y(n7),
	.B(WQ2_RPTR[1]),
	.A(W_PTR[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U16 (
	.Y(W_PTR[2]),
	.B(W_ADDRESS[2]),
	.A(W_PTR[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U17 (
	.Y(W_PTR[1]),
	.B(W_ADDRESS[2]),
	.A(W_ADDRESS[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U18 (
	.Y(W_PTR[0]),
	.B(W_ADDRESS[1]),
	.A(W_ADDRESS[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U19 (
	.Y(n12),
	.B(n1),
	.A(W_ADDRESS[1]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_RD_ADDRESS_BITS3_test_1 (
	R_CLK, 
	R_RST, 
	RINC, 
	RQ2_WPTR, 
	R_EMPTY, 
	R_ADDRESS, 
	R_PTR, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input R_CLK;
   input R_RST;
   input RINC;
   input [3:0] RQ2_WPTR;
   output R_EMPTY;
   output [2:0] R_ADDRESS;
   output [3:0] R_PTR;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;

   // Module instantiations
   SDFFRX1M \add_ptrr_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(R_RST),
	.QN(n6),
	.Q(R_ADDRESS[0]),
	.D(n19),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \add_ptrr_reg[3]  (
	.SI(R_ADDRESS[2]),
	.SE(test_se),
	.RN(R_RST),
	.Q(R_PTR[3]),
	.D(n16),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \add_ptrr_reg[2]  (
	.SI(R_ADDRESS[1]),
	.SE(test_se),
	.RN(R_RST),
	.Q(R_ADDRESS[2]),
	.D(n17),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \add_ptrr_reg[1]  (
	.SI(R_ADDRESS[0]),
	.SE(test_se),
	.RN(R_RST),
	.Q(R_ADDRESS[1]),
	.D(n18),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U8 (
	.Y(n12),
	.B(RQ2_WPTR[1]),
	.A(R_PTR[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U9 (
	.Y(R_PTR[0]),
	.B(R_ADDRESS[1]),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U10 (
	.Y(n9),
	.B(n6),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U11 (
	.Y(n17),
	.B(n8),
	.A(R_ADDRESS[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U12 (
	.Y(n16),
	.B(n7),
	.A(R_PTR[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U13 (
	.Y(n7),
	.B(R_ADDRESS[2]),
	.AN(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U14 (
	.Y(R_EMPTY),
	.D(n15),
	.C(n14),
	.B(n13),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U15 (
	.Y(n14),
	.B(RQ2_WPTR[3]),
	.A(R_PTR[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U16 (
	.Y(n15),
	.B(RQ2_WPTR[2]),
	.A(R_PTR[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U17 (
	.Y(n13),
	.B(RQ2_WPTR[0]),
	.A(R_PTR[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U18 (
	.Y(n8),
	.B(R_ADDRESS[1]),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U19 (
	.Y(n10),
	.B(R_EMPTY),
	.A(RINC), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U20 (
	.Y(R_PTR[1]),
	.B(R_ADDRESS[2]),
	.A(R_ADDRESS[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U21 (
	.Y(R_PTR[2]),
	.B(R_ADDRESS[2]),
	.A(R_PTR[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U22 (
	.Y(n18),
	.B(n9),
	.A(R_ADDRESS[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U23 (
	.Y(n19),
	.B(n10),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DF_SYNC_ADDRESS_BITS3_test_1 (
	W_CLK, 
	W_RST, 
	R_CLK, 
	R_RST, 
	W_PTR, 
	R_PTR, 
	RQ2_WPTR, 
	WQ2_RPTR, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN15_SE, 
	VDD, 
	VSS);
   input W_CLK;
   input W_RST;
   input R_CLK;
   input R_RST;
   input [3:0] W_PTR;
   input [3:0] R_PTR;
   output [3:0] RQ2_WPTR;
   output [3:0] WQ2_RPTR;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN15_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [3:0] W_SYNC;
   wire [3:0] R_SYNC;

   assign test_so = W_SYNC[3] ;

   // Module instantiations
   SDFFRQX2M \WQ2_RPTR_reg[1]  (
	.SI(WQ2_RPTR[0]),
	.SE(test_se),
	.RN(W_RST),
	.Q(WQ2_RPTR[1]),
	.D(W_SYNC[1]),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \WQ2_RPTR_reg[0]  (
	.SI(R_SYNC[3]),
	.SE(test_se),
	.RN(W_RST),
	.Q(WQ2_RPTR[0]),
	.D(W_SYNC[0]),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RQ2_WPTR_reg[3]  (
	.SI(RQ2_WPTR[2]),
	.SE(test_se),
	.RN(R_RST),
	.Q(RQ2_WPTR[3]),
	.D(R_SYNC[3]),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RQ2_WPTR_reg[2]  (
	.SI(RQ2_WPTR[1]),
	.SE(test_se),
	.RN(R_RST),
	.Q(RQ2_WPTR[2]),
	.D(R_SYNC[2]),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RQ2_WPTR_reg[1]  (
	.SI(RQ2_WPTR[0]),
	.SE(test_se),
	.RN(R_RST),
	.Q(RQ2_WPTR[1]),
	.D(R_SYNC[1]),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RQ2_WPTR_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(R_RST),
	.Q(RQ2_WPTR[0]),
	.D(R_SYNC[0]),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \WQ2_RPTR_reg[3]  (
	.SI(WQ2_RPTR[2]),
	.SE(FE_OFN15_SE),
	.RN(W_RST),
	.Q(WQ2_RPTR[3]),
	.D(W_SYNC[3]),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \WQ2_RPTR_reg[2]  (
	.SI(WQ2_RPTR[1]),
	.SE(FE_OFN15_SE),
	.RN(W_RST),
	.Q(WQ2_RPTR[2]),
	.D(W_SYNC[2]),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \W_SYNC_reg[2]  (
	.SI(W_SYNC[1]),
	.SE(test_se),
	.RN(W_RST),
	.Q(W_SYNC[2]),
	.D(R_PTR[2]),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \W_SYNC_reg[1]  (
	.SI(W_SYNC[0]),
	.SE(test_se),
	.RN(W_RST),
	.Q(W_SYNC[1]),
	.D(R_PTR[1]),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \W_SYNC_reg[0]  (
	.SI(WQ2_RPTR[3]),
	.SE(test_se),
	.RN(W_RST),
	.Q(W_SYNC[0]),
	.D(R_PTR[0]),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R_SYNC_reg[3]  (
	.SI(R_SYNC[2]),
	.SE(test_se),
	.RN(R_RST),
	.Q(R_SYNC[3]),
	.D(W_PTR[3]),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R_SYNC_reg[2]  (
	.SI(R_SYNC[1]),
	.SE(test_se),
	.RN(R_RST),
	.Q(R_SYNC[2]),
	.D(W_PTR[2]),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R_SYNC_reg[1]  (
	.SI(R_SYNC[0]),
	.SE(test_se),
	.RN(R_RST),
	.Q(R_SYNC[1]),
	.D(W_PTR[1]),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R_SYNC_reg[0]  (
	.SI(RQ2_WPTR[3]),
	.SE(test_se),
	.RN(R_RST),
	.Q(R_SYNC[0]),
	.D(W_PTR[0]),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \W_SYNC_reg[3]  (
	.SI(W_SYNC[2]),
	.SE(FE_OFN15_SE),
	.RN(W_RST),
	.Q(W_SYNC[3]),
	.D(R_PTR[3]),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SYSTEM_TOP (
	REF_CLK, 
	UART_CLK, 
	RST, 
	test_mode, 
	scan_clock, 
	scan_reset, 
	SI, 
	SE, 
	RX_IN, 
	Tx_OUT, 
	Parity_error, 
	Stop_error, 
	SO, 
	VDD, 
	VSS);
   input REF_CLK;
   input UART_CLK;
   input RST;
   input test_mode;
   input scan_clock;
   input scan_reset;
   input SI;
   input SE;
   input RX_IN;
   output Tx_OUT;
   output Parity_error;
   output Stop_error;
   output SO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire REF_CLK__L2_N0;
   wire REF_CLK__L1_N0;
   wire scanclkref__L7_N1;
   wire scanclkref__L7_N0;
   wire scanclkref__L6_N0;
   wire scanclkref__L5_N0;
   wire scanclkref__L4_N1;
   wire scanclkref__L4_N0;
   wire scanclkref__L3_N0;
   wire scanclkref__L2_N1;
   wire scanclkref__L2_N0;
   wire scanclkref__L1_N0;
   wire FE_OFN3_scanclkref__L2_N0;
   wire FE_OFN3_scanclkref__L1_N0;
   wire FE_OFN4_scanclkref__L3_N0;
   wire FE_OFN4_scanclkref__L2_N0;
   wire FE_OFN4_scanclkref__L1_N0;
   wire FE_OFN5_scanclkref__L2_N0;
   wire FE_OFN5_scanclkref__L1_N0;
   wire UART_CLK__L2_N0;
   wire UART_CLK__L1_N0;
   wire scanclkuart__L6_N0;
   wire scanclkuart__L5_N0;
   wire scanclkuart__L4_N1;
   wire scanclkuart__L4_N0;
   wire scanclkuart__L3_N0;
   wire scanclkuart__L2_N0;
   wire scanclkuart__L1_N0;
   wire n12__Exclude_0_NET;
   wire scanclkuarttx__L1_N0;
   wire n13__Exclude_0_NET;
   wire scanclkuartrx__L1_N0;
   wire FE_OFN14_SE;
   wire FE_OFN13_SE;
   wire FE_OFN12_SE;
   wire FE_OFN11_SE;
   wire FE_OFN5_scanclkref;
   wire FE_OFN4_scanclkref;
   wire FE_OFN3_scanclkref;
   wire FE_OFN1_scanrst2;
   wire FE_OFN0_scanrst1;
   wire scanclkuart;
   wire TX_CLK;
   wire scanclkuarttx;
   wire RX_CLK;
   wire scanclkuartrx;
   wire scanclkref;
   wire scanrst;
   wire RST_SYNC_1;
   wire scanrst1;
   wire RST_SYNC_2;
   wire scanrst2;
   wire _0_net_;
   wire ALU_CLK;
   wire CLK_GATE_EN;
   wire PULSE_GEN;
   wire RINC;
   wire DATA_VALID;
   wire pulse_gen;
   wire R_EMPTY;
   wire W_FULL;
   wire R_DATA_VALID;
   wire ALU_OUT_VALID;
   wire WINC;
   wire W_REG_EN;
   wire R_REG_EN;
   wire ALU_EN;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire [7:0] UART_CONFIG;
   wire [7:0] DIV_RATIO;
   wire [7:0] REG3;
   wire [7:0] P_DATA;
   wire [7:0] SYNC_BUS;
   wire [7:0] R_DATA;
   wire [7:0] R_REG_DATA;
   wire [15:0] ALU_OUT;
   wire [7:0] W_DATA;
   wire [7:0] W_REG_DATA;
   wire [3:0] REG_ADDRESS;
   wire [3:0] ALU_FUNC;
   wire [7:0] REG0;
   wire [7:0] REG1;
   wire SYNOPSYS_UNCONNECTED__0;
   wire SYNOPSYS_UNCONNECTED__1;
   wire SYNOPSYS_UNCONNECTED__2;
   wire SYNOPSYS_UNCONNECTED__3;

   assign SO = Stop_error ;
endmodule

